XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����q���(�äɶ�����z҅�s�K�h�ʓ���=R�o<7&ɻ����B5` ��ͬy��{���<ĒAx
���F-u�D\aL c0���$�%�:�?��Ñ_�ը�+�BsU�޵*@�� ��s�N\��
�/�l�WQ媶=����C5�gƫ��nʹ~:x_E�#�������Td��ûd]1��3����S��\>�L>��w0�>�;W��+i]�Ѥ�؟���? �'��/8f�(zK Ђ���Ć9&�v��~�Z^C�o�3�II{O�O����-T~brޤ���6��&�o��9��*��"�FfS��Kon��)a8�A�n���cG{��*�@�Je4�j5T��m/�A�ЧX"-��x�̉9'&4�29J�+�.A��L�(_�4thm�-&?�>i���%'�"X% z�%=���YH@eρ�ADr:��^\lXQ2�P��K��?YM�s�H���_./��g�-x������%�:�o��e��8�x�����\��nfT{{�O�vZ@�sK\!�-�����V_��}d�a�_/�)"��Y�ü,�f ��ǇJ�Ό�ffk�h�'��R0.q���q��.c�	g� �Mͅ�����!/���LP7;�kp��E������C�K��0��x�!���ab���~�E/#ޒη1/>#��Π���^ܸ��a��S�����B6������Oמ0W�m0�q�A^o�Wp�TӇ��4kr:z�l���\{XlxVHYEB    b380    1930����D��Ph\�1
VAH87K�|p��W+hڳ�ʝʼL��W��ל��[��'�����(3cH�������S��D�L��6�K��h?�n�.(�/<�iO������)_4˶�3ea���[`�	l���!!�S��C)�︮Y,})��J�^&���m��P	���0�Y����^���#�ê�T�l^�� ���u�9���"%��	P7��"mI��I�]�.��zݢ{��w��`/�8qL`�t��q�_������ֽ�0_�<P��:�/|�D��Jj�O�h���,<������Q1����si�&��t^���q��>[��s�������M�]86���!�r�M�}1����7��*�#��[I�(Y�2C2��mg�7I^�B��n��#�G��Z��2��|.hpv��60A���7������d��o���
���{T���[��U'>�5��UϪ}ٵYR9��N���]j�<��G�/�e�,Km �~��㻟E�b��4T�:���V������>����Rk�0�&m����J�-�j�IP?�!Y�"�q�.ܢ���5�q�"]<&�֐�ڊ=sO��#F_eB�0���l�'�=iXeJ>A�>��"(!���fm#�{.޷�7����M����a`N08���mv{�Oy� qrp�O�A��j�1�J`>�ʉ��xl{C���ik0<���t:��F��������|+�;,װ潰b2�/��m�Oc��&9��j������$zU@�N��2':D�G�{���X����}1S0ă��Q���w�e�!Co����`����> %���L�h���АN�p]ɸV{��g�;l��%�vvuC�ݲ�ֵ~�u���4�UR� �����X�t����-�_W�[�+N��b���?����8�ě�%�֙j,4,��I��3��b*����z�Ѥ)�������.��a�i2�A?Or�)�gw���;��R����ؤ5��w����9�
;��h��3í"�1?#��C�R:����D<dV%3G��ćB0�5	`Y���v�I`nᔍ<ҧ��Eg�4�~�jp��X.������5�	r��8)ĸ����u鑋� +��$�b4�ۄG�� :˷�>2*՞���+𱚮;:~�eP�5�����ǯ�]0�D��R�>��2|@?Ͷ�~�8àWO9Sl�7�'G�sp���
�)5$��Ss�)�g�myZx\>V>�|�t8h�p���"<��XK��h�=��Y��Q��LT>P�ǔ64twp���[��[DX^��(��~��
�Z	@?O_*���ȼ�.�d2e����Vr*`&���BY
�My'@]��%ؼ\K�vY�	��L�ߠ*S7[����@M.$�9{P�E0ĸ�.�750��n��>��Q����[GN�o� �e����Һ���?mL�90_��v[��P�b�+կ)�G�I�z��VhN�*�~�������͠A�x�TDJP�W���S�.9�}Z�Y'ا�՛�r}% L�&�
�o�=ɔ
hk
4<�H9�D.%���OE�S�,~!�Or�\4�^�Sh2�v�[�\��������17έY�Zӧ}�8�+��OA�<A�(-8�!�,�}}��P�/�_��c��X��@�(�c*��Z���S@y�������B)[�^���~ZH�T�~{C=�����y��WY��xf��n]!��n�������B9֍Bn/{�l���6,/�	��f84�u�k�����0�F�e������W�cf�#@�mk��2�\�D,��c:���\���	�t5��|�$N�9X�bC{�kw�O~�Q�3�>sm:�-�����9��˳�V��������&�pv�ޢ2�p�T�Iu�iUg��� �GZͻ�S-ߵ�_L%/Q�hx�������묫*�o�q:�7~���+����g-�7Fn���s\�jߍ'5�^�Ԭ�G�����r_t�~a���탃�	�7���H8A�P�C�$�wn��*=+d��b�t#v�q=j��w/X7Md|^�Te.�s�@�(z�
o�v�����*�+T=	t�4܊S2����Pк�1�3KѢ4L�;���&��Y��O���T�8:Z�,Z�W��&CC�������F�X_��k �:K�3�A ޫ �]5�q}:�H���x�wAX0ܒw�-��q�L�WM�)�^���7{\hZ����F�Љ��8t �'9�}X�m��X��g��;� �p]�
�ꖛ �f��D�ź~̸�MeD��v/�p~�jeY;B-�f�[7_ق*�:!���	0�����ZSڜ���I;����}�us�-��$�3^��U�{_�+��{�|�>�Oנj��Q���y�<��A��O�8��f�
Rţ���*�b�t�c/��w��O������ ��G"���MLi�y�6!���!�Y��t���Lo���N!9����]
H�$���U}�=�4EYY�ʆ��f.*tL�}Js]�~��*� dɌXV8g�r����!0�P�蚋���V�w�o��b����g�Ƿ��	�q����$�Ut�����}LoSa����T�~�^m��2AS��#�/l!v�W���?�7�i*H\�Vu�r���đx??S ���Ӝ�Q��s�:�]ݔI:Ð���2:6�gpEAV��6YH54�V2˳��R���e��T4��˖���_�KK|�,�z�����!w��(=s��0b��W����	�1�_��ݵW\��� ���h	f�23/�雦� �?�(��dύ?��>�KF�.�����C��yv\L�H`l��ߓ���mq���
ǭ���:Ͳ��Q���)b�NQH��:�Es�A�^�>Hu���6%I|H�ҐPE��0���9�����H��JMIM5�Y��&A��	�N�T$1�w�V�6w<)0����� A	��@y�n���Q��Dʏ�'f6��wʿ
A�H�.���T��Ĕb|���� `������q/wBS͌���f���� �(����{,u���)�D��C�핢��&.Bi/t�^	�&������
Xu���Ֆn��sظAF�N�ӎ�6� �f��ld:�<.�{-�?��\	(kP�E���u���L�5����մ�O��Z���Q���z����6SO֍��ԝ�G�Ł� _�_b��X&�y��!�^�?����X�8�<���m#q��"*B�M�dr;@5�n��/����t�pLkI��(F�`>���d��*�ު�/Dʘ�l�s��؟\���[����ey�ȑ*MU4o�^���P|#𾺟�8�r��x�+���.��l���b&�g$� ��?��_o��+c�n�&�h}��x}P?�eF�U:��/��5=)���,���W f�"	���i���Y,J��Ƕ�ץ�&��Aq���B��Z|���\�,��	̪1���S�e�IPy��d�?�2�&k�`���&�;����:�%�XN��z��r��^�9��S4��
�<��|��of�E�yr&��^ڮ2�7C��ˠ�3{�>c�t;���7�)������HZ��y��.�����t�W�����3QmRAxF��d��7oq�gJNz�f�{�5�W�u�?�o6|^��-����M:]�W�{���m�8n� �a�C���a��"�f�Ez 8�^ڑ�J����`�ѓݣ1�C�Ƨ��!W�� ��=�K��:r��#�;l69��sd�{,�����R&���*!�!�C�/�"u��i�4�N�x���{�fPk��ܡ�y���n7 �1Ua���I��ӕ'0@�O͔�$�s��w��w��=�@�X'��+.uu�jv$����	�gc+��a��uPP�1�& ���C"�������KΖG�)Oi�8���d��,�dX �E���(4N3�NcgL��+҆�>�l�Y�Xh�D|&�k�Ė7�
Q���z]?%"=S�e��;p�wvK7�$L��ir��Vf��x��qƸ�0��мւ�n=�g����]���)�RI�!,����y�칎e��sjU�I�hO�)����1T��V�_�l:�iU�,
+�]7���(�E��1��|��L��[���t"&��(�����m&P ��oa@�l�]v7�2F�k$q�S��ƃ�vb�e�F�D�B���%��F��/��:鈶��ھ��-72��~� �lp�s�ӯ�Z�l��P�=1�3��k�t���_�Ff/�.�w��1K�7����Z���#���Ą'N�A4�
��R�}g�f��P�5v`6��*�c:�L�<ɐ�x�@F������z}h�[WE���wL�wN7��@��9EdE(S�6�2��$%m}�9�d#�7�b9�W;�#��������Yh�y_����.���|Ee��q�΍�~�_��[���w����V�5����K���%�z�"KV�_nBߊ]4s����n���.��g˱M�i�st���
e���FO	>��h�f�7�>�$��-!,�r�X)<!��t4#�#�W�W�
6�ub��i�e��9�Z�ÑOֵ��xmx��6�gщOspѶ-yLK�B�p�O~(�V�F����-���֛�Q��L�f)?��"���&��D��GE�)K�?C�e�c˒�hwIB�*��󏞕���;����\�.Kn�ߔ�ua<R2HN|��N��6�5)�,d�-������(H�{B� b�=��<~�VN5P�����gr�w~'���W��n��| u��o��+�G�sc/���"��h#��C�܊�J�'�¤	�ѕ�l�nY�dC�.V`?&��~�?U4`ƩU��<�?Ҹ3�V2��F�e�']&h��(�y���F��\�K�S<����sSXE*���G�k6{j}���ʴ��Wl�?n�,�|Kѣg�h0�1gw���`t/��/�/1^�}I������!C�"e|��9h&�\)T�<ْ�m����P�Շ�6v31c�i��7��������'�o�Q*O>C>K%|u�0�jt��|^}�S[���5�������T��k�;[�۴���Tdh�_V�m�;v���%�Y�J@�9� �	�������A���X5�3ڊb:����tf} �L��vQ���%1���y�3+k�!'�dm���L/�^
6]�E�-NLa�J�6���2�R(P_-D�C��|��hHF!�0ml�"�W�?��M�]��O�֞D��P��X�D�'��;)duK <����p�,�No���Y(NW�u!j��
h���\ۭ�[��P�uA,/;�u���m�+�[^y\_�쟙�����S� ǧӽ~o�G
=.W�o{ͭ��Ҷ�X�y���A'���E�Y�S�6�X�詧�����3��ʧ�ǔ����V�8�x"�����ƛ�������x8+���V�#�J���	�H�wn[�ƀ%��m�'������_p16�)e�
��J������+��%��C)�M3%��@|���[�:���)�;a�ȁYZ (+���L���s��q�t(����X�:�xy]�	�tۜ1(T<��x�x�Jf��(W꬇�G-(�Kdk�=�X���� QX���/WŴ<�E�js!�m�z�6:i�����K���I�Bf{��>��w�Mu*�j} ��^�$}ar��%��Q�ݿ&�����}}��"��9RF�VY�eh|w��;�#}?$gyT�wi-[�zQ�Q���m��-tw�R���1���e���Bۗ�o���±�@��]9�n�HLXuV �ϖ�w����c�k�GG�h���X?�5��4Xx�@o>����`F��$:�b����2_��n��3��@�&z:�%!�j����ڵ��G�/	z+y��Hr��w_M��}dl��d�\ ��j���?JT�&�m� $N<g�՚U�����ݘ]ƭIBh�<V�ջ/E�����H�����Zb��=ܥ��E�HI%|��SAK�)��I��$.U���*��T)�:�\T̙r�A������E��$Ϫ8̕hуb���+�e���|��W�L����i�	��3[߃����������.�oI;�>|����9ְ�z0��e�����dM2+�x#�s$���o�9�*��d7�5 |��_�[�܈�RcT�ib�9�]n�8�5�
x�� �s�u	[�:{ny:3�i�^O�隯D툺��v�&�r��$����H�o�]w��W<<�H��Y�)鞸B��5�ܢ^�^��/�^)������k��&�[,=+"�IK