XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��7�R�r�T��#! 4(E�LP!���������Z>���"�C��҅2�6���_�����O��\�/��/��B㵄��Q�'x��p�B�`��/�iW��Ѷ�么3`^�Ǜ�b#�,y�'&C�����	1fL��y!li�~�*�QL��`�s�-�C�ܦ?�gU?�t՞����"5�⤋}�͇��������ǰ�������ۘH�!��Op �Ae����+;�Qh|:��{�-�c�p�uy��/]��d�s�O�<�����a�҅��*1w
��ӍMu �Q�	_*8"���z�Ş$�g2�<ϰ9Hi�����y������k}8]���\f{��.�=C�� c�P�t�<� ����,��4 �t���bL)l*��0[s@V�:�j0���c4��*��	iǞH(M�O�<S!��7v�D9���q�ޱ�!��Z�"��Q�f�p�D��MP��0��_����*d4�-#����ֻ��ӄ�;�������c���7��uh���"�z�;����q*�t��q��
+��H����rǋ2���y�a��%D���1+���S$&B���r�f�@�'0�*|��	]ʆO�C#U!+Ճ ��ݏ���:ݮ0�:��ꩤ��܂�`C���ݯ��I�����n��"mZDk:>�a���F��$�^^�X;��.�ߋ�����ܘ�G`�����}h��/�LB�Ϋ=�y�B�Z��3d#V���U��͸��`�CH2�VO�8��XlxVHYEB    33bb     c90�v��E;	͠�{z#��H��f
4Xh��S�|�<@����՝Bj�E��="��� �Z`�pZ�c}�tN���/�On}&�]5��t�L�ÉSF�j/���A�rYF_t�u�7M�Y�)R���1g���63KN�hx�&���c-(dK���!��0״����:� l���<�J�ɏ��Xjt�Q��8�Q�H{���'����G䷍�8
���2�KOE��a7�d� ��	����OE�䴕�)?�sV�d��'J{(�B6x[(%����?O/JQ����°\����=v���G��7��x�@q1�Y�lտ(������h�zV���@[P���#�棱�s��7��{�v��z������B���$��<�� ��GhqWd�B9*�����p̚��9
4�@�G��S�X���Viy�ʴ�=O��v�D/N5B+_J����᥎��� bH����j͜Йp:���w$�蕵��1����4�V)��#�L	Z� �X"�꩔�TK�c�);>���aic���͟_A'�����#�P�\bz<È� ������Ӕ ��1ӈR���|	�4�	(v���E���oٴ�H ���gi$ropG�B4�����@j��Rz�!ʎ�+6%�����t�/d����)��2�V�j�)��#f��̪a�O��]�&��g+7�g�E&D�}�x�He�A$��ʐ�8�p���'i`�mp/��>-��a[�NXj�U�jt�f˛� ��'���1q* �Z�.��4��.�b�K@�E�<�Yʂ��Z�!yF���V�����Q�Yqa��"��U(O��0� [ƶi9�l~J�-�䷥L(cN*S�`�d��[��,�hT$�%k��K��U8����2j��.� �ֹi�����B��z�r��)>h���J줸V���%�T�yM�u��##'۞��
�=#d�a;/��Y!�s���{�U��;�F�&α��.\�֧�+�QD����=�;����~�֭���� ��jd����Z��i�VG�W4�&��h�qɄ>Ȥ�#�~p��f����3D��U�!�6�� ���K�-B"��������(Lb�,}�q(G��a2sJ�#�'�x�m����-w��'�p����u�D��ʍ#%�+��B"����F|3�?/�[��~k�+�x�50 �0�����t�i�/^$���e���zn(_�=8�	��a~#����U.	��
����f]�vb/%g�7Q�t�$u#�HGC���;�gQ#t�q8Ԇ����{F���"@\��)8��U.�jv/�燐k�!��Qz�͆�pǓ� �نA�2s�x�^��(9:M��,+����:��8��>�J1l8(z�~ <N��-��_9���J��S&��Pdl��>1]
r�(?�N��]��ڝ
V��i�MI)�"axx��*?�yŽs�O� �$����X��U֙a�o�V��%��6D%p�p�1���$0s�Vd4�	y�FiO��p��uW�D����O��S��+q��$�b��8l����Oʾh��:4����6�G7h����I41[�3��k��ܖ�w5o���@<����}�6����mb(��4O�y�3,S��9a����ז�"Ǭ��?��XQ.����"�m���Ĩ��<��(:�&��e§�(\��g����8��z�/��6���VAXZ�B=�6K�$���zaE �y�j���N�\/�b
�/��U�t!�Z���]�$ne3�e���,��r~q-�뢣�����v��d`/�
BF޸Z��(�"hC��=y��=����,������8�d>�!�E�Q[E���^��1$�6��!23����� �~����u��Izsg���mQ��9�&|頥���k�t�#���z�~3���dS���o���KQ�C���*zz�}��"��ɟ�fE�2�}�$�$'�����Jв�}e�I��pl0��G���\�K��K�^.���@����&�u'�|�1L� ��:ίEt���61��)����؍9^C7�$��79C�u+�u�DwLb�&�k2ܖO�N��H"�nʊc�0J����+7%p�����m��0��Q>�XI;1��x���UI����������B���{�1:��˔Ի��p1�.�yL�K�5�LS���Z5v�:l�����`�" �{ߡ�M
l�D�����+�8�צ�K܍l\�"����c��L���LH�Sv��wdz���_Z0�H��Ѡڛ׀_��Ի-�'��>���+ɡ�y1�!�TZ����C���(�V�
�����Pie��L���2-p� �Y��W��B� K�s�g &�G�8����b4s��g�����ul���Q1,�\wd?���ӋyV����NO�pD��Xyw�7�>�6��S
�no�Fu��QA�/�.�X��>�?P��y��< ���� *�����#!ā�޿l��<2um��D1�3��ʸ"}UJ7�����Z{{��tU�|���	7��h>m��a/Bܸ�(��Zz�@�,L�$��������������ӃP�;%MiG��ʊ~��SB<�j�n�]�yw��I�.����$��x�@��E�2���Y$�mkM�!b��x�/����c�o�b/���S�%��ʻT����Wޱ8 r���\�5>�xb���8��w���=g���?T�L���Y6\�N�E�^k�n%��ġ*)f��e�#%�a�M�[N���x��s(8j1�X�/�T�g��+G�,K��Q���WJ_�&�z��F�2S�ǋ�I�)l�،+I��������f�2 s��c��@��+h{Q���Hv�}�y����ecM��n��N)*�7�s��1Zo����8�[���a�N1@�x��������"'v40�hr��e����d�H��x� �|�Dl��bhlB0�fg	���U�R��C?-�N�j�:#�ɥ3��_���C�k�.�����mM������7��\A�O�{��K(�ZH����.��/a�d �3%�5-�0';E�4^Q��胓h���J�1�o��RFn��o��V�O0��sZ���.Us�Ӛ�T�^�c�Y������W$����q�k Sk�}�7X�