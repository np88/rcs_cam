XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��=��j�Q�2C�3^�H���i�6��C���h��{�`�i�U��$ꍚ}�Y��j��N��8Ԡ��]K�*l�	�^�נ{y[��,ߖ*�RA"+4�L��)����ʆF� 7C�C��L6ar��� [�Qz�W��
B� )6��:��I5��d�G��O�eJYt�Ϡ=�%ȥ��8�F]#HΜ�Q��/�%���_���]mG����aX&c����<C���7)Z���I�pu�N�]��FpGp�0�2�dzd�x7�J�q�b*��������ޥ.�!�+a+���E�q]��1���3 Q
�R#8��$�|kG�c��[����I�����'�O4�4\o��	��-����lVܝ���(�7ۮ��UzRMo�O/�h�e���t����C{��n�ig����Y�nkVӼ�Z'z/ߙ���Y�;\���DS�z'�U̱~���"3�� ��J]D��aU���Yg��\ɗ���]�|Uz (tW�� )��,@��,zG�HEE���%��a���(1���Er�����^B��l��C����-O�g�3����1;�/������}�����c�b�=�0A�l�"���ίQ->�����p)G���Z�/|��pz�c�$����C���(���Ⱦ�ڀ�&���������B��6�������W;��T��.�N?���v�aϴ<#��b���s�yT������|L	fF���&����F5~'XĎ�uH�$�����9�3�����myx��XlxVHYEB    25db     b60mU����}.;�2Ⱥ��oj�lj#���%\�������tA8��M�#[�"�$�wH\����;l�����a�ZI���a�U��.�U��X�3B�a嗙x�i����3�+���2�$~`2�lu�Ao�#Q��9ӹ+�p��%Rz�
�bY��/t�^��C�������5M�gTe�0�F�������'�d�+��ٍ:$�k8�s���5V��CڝCA�g�>���]�������PD����j� �dnx)��j��fWYG�'q��A�����6�B"�\/��E�����49΢�A�DK�s#�;l� ����D��8�	ME��9�� >Ͻ��|c�[IOx6��=���{�*#�!R�	�gp�mGɝ?��#j�g�M��N5������ (�r�3p~M}�M�O��W���� xv�Y}ȱJ�~\{M��F�Ӏ�0�L�\�%�zv@A�0�?Ul�X$�0�_���r�Y(�E�L�?&�/<�oF5�e�d�K�a8^�R'֞������0��C?OV+���Z��v�5�����x���6�uI"�1�-~����a91�mW�o'�ȥ��ڈE�7e�Q��H�qإd0�H�h����IR�u��+/��9a��_UЩLg��ڮ����Q�R���O8ONi�o,�"����v��<��M�pAD��B�1���3��|�R������U�����nY���li��ձ�~8���P�� Mc8���i[:q�kD�œJ�����D`�骘��.L��E)��(��2/�bہ�&R��A�WK��9(�s�SBkq#�?���AL!ty{v��?V�51�Jcl �:d�)�g��%s�_�{ﵙ�M +dM�Խ�iy�����!f�� �Ej	�n�j�k�ʾR����z�Mߖ�x��yj4���8̂e~[��  Q��n�*�k��l�T����빯�V�~r�Gձ/f���^��Z��R�4�! ��;�3K,����
�"�\_n/�HG� �?�}/��#�oi�ݿ�:��ן��TU䱋���1����$�'ϊ��0���.o�s
fm��Wvk�X5��Ux�O�o�������H�4�/Xy�^p�(��']�߮��i�1-�ᱫ��}�x2E���r�)
�5{;�4d�]�H�IL�5���MW���S�/����~`��ȓ���X͞kN����O"�����4=�����r�==aq��\�wȳ�%�x�R��L��Iz�~v�H[U��l|�D�_�Wx+I�-�*E ��YPOb�K�n?'[8p�$j䓲�ɟ�������w>`��G{�=~��T�O]6�T�D��m���@�,�3���kښ�ڗy0Xn.
���u��w��N�Ym�+��a��{�ʄ%��� "ܬ�psf��û�1��v��P����_�cߡ��V|97�uۤ`͢H�}���x�B�|"�8V��d%�b�eHdl�rIf�Ψ\���6,�ǰWxc$�P�kF����Y�o+��tv;EX!JdQ�2&��M-W�5�B�8�B��fv`:��y���g�
>pq�f[�˄�A��Q�=��<E�9���P�Z��r�F؝{��P]�
�=s���7�[���q��>f5J�15ר*]Л�,*#�FM�du?�U;��1��Q@;��ϖ�o19S2O(�Y3�k�s���M5�2tHƔܱъ��Ŧ��Ɯh\oRד���$�TH6�C� �ZQ��@����7/2���|�6��
;j���n��1�$��H�%g�p㇜ϝ<�4��i�ͭE���+�u�^������Hf�i��3��v�UY`�/��`�*��\V�<����s��G �&��{�0R�D^Y������1�9Η�&q�heP��)l�bFj5f��w2������g<����X�Aж���φ��b��s�'����<Ș:�Z����q;�CO�0G�E|�<<.�,H�����)��c� �J�9AJ�T�[]���%lX���s����
���lm`���N��f5�33��k������Ԉ�Ms�Q�:jNP�#�0�҆�Z�V�3�OL߲�E�6�e�qG=�e�����J{�¾��c�P���ի�E��\JC�������D���;H�@�=�ނBr�
&��2.��[��`�D�o��	�FZ�m�ud�K�ݔN|�{%(��"'�z�2Ĵ��B}���7r�Y0��f����9�o67�6�g8,��ﾐR�v�z��ŵ��*�lͯX:����7��-HG!���̶�R�ӧw�.%�mpHW�}���mh��&��dA�C*��ڦ�Y��51��/��WN�s̍��B�P��/�xi5�4j�'�-5��u��b��?l#���A����Q�,`ND�TѴ�Ɓ������u0�`(�i�J�� !%O��
�"�*8R^PK���q�qx�a7^C�ݡN�`Y��gJx̖	���.ma����L��B+�{���K�,7|�	8�+�u@�ԇ�E�`�l�Hy�����4�^f���������|�NT��y�v\
Iע/�G{�+P-��B�qk�P�y>���p���4��+�@�;ՀC<�
��6/�Ԣ��n�*�� ch}E ������ąQ����IEǠe���]��3�XU���t')���D7]P�qbV�r?�b�o�U�b<�;�sE���ǣi����tM����-���+(�|�e��}z$�Ԯ��	�2iZ6Ya �~��3����!�����R�J�'���XKO1�܁/������UP��"�6�_-��B���ƾ+�\�+n��1�9��cn�b��o�� ��4�{LѼ?���&Oq�kH}|CQ�?�W�y