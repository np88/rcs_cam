XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����o��[ \_�'�%��K��lt�\������:`�^!�w�~Z�znSx�\�Ў��MJ��+��b ��l|�l�����D��],�!�����U,U��{E�t�sp����$�v;jA��
�}.����7�a0�D���]��嚪�^�	���)`
 �o�@��'\ݙ�r��)��aa�U��P��9����"�S�j��h�i ���F���B$V�N�+�,x���ր�Ƒ���-}�l��q=���-K=Gj�K�}n��E�
�`hd��3�m�������}W7����?������	�~�&��hϳs8����J�Б%�K69�D@�oI7�Ǘ�RI8���V1u�)*�kÙ4:�x�=�/#J�'ʂ��Wp@t��d6`�b����=�^���4�*E��rZZ�j�2ԥ�C��S*�����g�� �����]��/I�	$6ӥ� �gW�P���,�v^&��n��W���;�Lm�b�l`��+~���[>⢏��9Ѡ8H��;gp���b�9F��s6{Nf�- L�_�|4=��`v_��jdz��N���5�1�C�r�F���?5�ԛԔ��`┓��|A�ȥۦHШ�ߴxR��K�g��)uF8�;�_?b��W��`�����\�"���y�).2�s���J�a,��qu��/E�|�Y
�6�,��uK�a7���?f�����Kn�)�*��;�H��>�������5J�J�+��C�؍lt�h��u�XlxVHYEB    8388    17404U)$�/b4W��A�3w��ua?�I<�ڃ�s�5�Q��"��H{td�G�
'�#�[�}��M�p#�]sr,��#���E��ؙ�L$�Q��v����V�72Z1R(A�������Ӵ��M���p0�,��.�����A&{� Kʣ<w.DL"�o�+��1�����l6j����t�{3�yS���
LW=)=� �K�\������jBI����~w�g�n����dĕ= x����G=�r�U������~���!V�<�gOb׍�'U��!w�=	lO�J���V��FZ�6����'�7���Í�8<�ř���C�6��Nu�T ����T८Mr���ؠ� 7�Y}oto7��j(BV��
�� ]q啩
F]�+��C��E7��	.���Ff�\�=��N)�Ä|�_~�d�Q��,^j����V.UR�niL��T��o�ј�Bp�b.��gjxN]����y��
��Vth(By�s��T����X���
c'��D����Zj12u� ��^A�O�6K�g:#��O�
�[P�H���1�Z	n����A��R�T��V��(b����L�fa�t3U^��(+A�����.*;��U�[��������%F��D~
���&6��z�1��<@��o��P�(�m
*���R��Vբ��c��&���1mD��_���(�R�U9U�}P☥<
�8�B�����A+�!�ִ�1���+��)Cv�^���3�+p��vgq��p�f�՟>�?�`p�(;/N@��'���3�{���IE����<%͞�D�����|#2S���Ae�ܑϐ2�q�C��j�w�b��8���
�r��D��^lɏ���i���J�E���gh���p	�䯛bwS2�8蔖>c�+,�Pzr�%!#�a�=@h��8$iWD9(��`��M׮�*We{��[��V�M��QF��D�Z�#���ٮ���Y@�⊹�w�	�Q��U9z�ѵ�(/���R퐐�e+j���x�.́�_�d�)e�
���Z"R���ː�
s��ol
��H�h�'NgQ�/ʊ�bӌ�
{ٗ}_�t�#?[�_������i� �*`��誕��.�\o���5��Tq¨�MI���f#�l�ȷ�:q}�$��D�h�K��nzV6�� �&:��s��}�Z�M-�T��Q'i�5D`�ϯO��|��E��#2b�s�V��%K�o�Vc�����Y1��Jޕ�Z��nI�[>��i��p��@�<�y������ekSPˁZ�(oD�ʹ;^ٍؒ���|�~>c�kc*$��&<�ۖ�ν42�^8掤��.�/�RXi�-X�E1��#�M������g����4j��9�W���s�:Oz$�Y`�Y$�� ��7�V�PЂJ-~g;��ِm�_]S䱹)���OŔuCW�I*2䱷��Q��9�p@(9T��Rx��+�-��E�q
��M!�3Y�.�z0VvrWA(�]Ra|K�l�2�6%&_Ƿ1��Lim�]#��Y������]��w��#�#l5�ؒ��I�lK����L/0�UG2�H��&�`�P�}������1���D�E- vJYSz:vB�h�M�Pe�CaJ���������g�� ���V�a����P��H�CB�/�T9G`�Y�,6���F;&�2z�B���eR+����j�(��I=�J�+TN���It��8�(�z�D(�Wi�<ST)��$���H5=�?$���W�m�uT]g,�}Vt4+�d�Y��1{�)V����X}�άAS�".�[��p�-oR�`�H��!Hu\1Sj�Q���&˼�u~�jb�����Xs44�'���N!�!%��p�����ݍ��ޕ7+�Xy�bN�~[��k�=�|;��� &�*�����_(٠cC�h�N^ɗg���e[,B�e7�3�弗�[�0��v�G� 5�@!�ca���K�/{c-��O�æ`P�
>i*	�hu,���˷U^�z��{��f>�����޶<決�~��ZgD�"Y�6�A79;�YḬ��D#`b�7d�bA'�j��
�����6��(�W�=�X)�IE��w���Ml��geOᘾ7��hX9�11���M9o��F�Na1���@+�� ��Dߟ�f�,�c�FQ������0���s�fPHSI<�&	e���m�X�/�oٮ��_W=:���ij���0H*��߼��l^;-r����M���[;3�h�j�b�
<e�EZ-Q��ބ��	}�Y����1�uM�������͜�|�n8H���T��Ⱥ����6�d_>(��i9�[�{Oّz���T�tJ��b���o�T��͜�C��rԌ;P!�\��5+�N�x>���p�2p��������
x�{�n�����U��2s$��9��Dn5��+j�Ƣ,r5�?���=��I�4���r�����1�00K���'(g��{m����7�{>
GA�xL�Px�7�[e,�b���Y+���}��/����ⴆ�w��cW��! =�d�'L���zlӡ�tv���$6RVȔ�F�]h�T[��F�x/�Vx�'��h�&>�TF��|�i��.R[�W�PUzY���]pX�T����9H^+r�M���lJ���9Ζ랢�ر͈�k���KQQ���dM��9ps!��B~��5KuZz(Vϝ����D�7��U~L5��;E&�C�4��g���2�|������0�C�Qֶ��~\������R ����E�M&]��6X�ׯ�6X]�1J��b�Pd�h�P�M�Rͭ y-ˉ/���R�[����=`����Z�`t�����9z�!��н T�-�0)rX�Fdm2���$�&:��x.�ך�Z"�S�	ɵۢ.Z��6�[5�?�c�����KV�oШ��(� �F
��Z��W�מ��?��)��B��{��-#�����f)r��iU^B
�C� ������Z:��A7~q�$n��K���I(^����4wl�'9��ڣ��mr
8R7W_�ԡ������o~�i@4����'�i��E�WL�L*=<� ),�5,�5�-#(���4����EԘ"i<�3b��<a�D�[-_p�ǉ���~�0U��F�$�w����A�}{Agw�6���x��n���������L�xKN�x�fo')�tS^�^�L�]�j쿉&M���Ak���a<E!�k_��A���>]#��Ov�����k���H�9܀@��� �k�v�۞_��:��t$������R-w�0xE�$�-�ֿj?���z�G��B�^Ԅ���r�a�R�FC 0ۻ�E�z�5��DYŁ���&J��8�B,�_B_����[s^��x�$���%�v1C�귰n���V!M�q�yܹ��D���ݴ"�p������d��2i�_���������=�q@e �Z����;f�|�۾����c��J���F�Q��vuZ������זVcRS�QgL�ךgP*�Ye3��@S|�\W�X��3�a���<����C&�Zo�l� fv�����l䧓��
�d2M�衖���]�P5RQ�Q�w@}��{�V2�e��Dױ�� �e=y��g�����E>����:�g��a�5hJC��L{�]�S�XP�^&��9�;�~���r	t��(�d�X���W�(yS���.�ʈ�Τi�PnR��*a��5q�{�i]�jn��e���5����o<S��z�EzS��7��h����B�M'!�A�
��'S�2_r霰��\M�4k�c�b�q�z�v�:u������='Ⲣ�����`�24��⫘��,��,��(ڬø s�Q�\���ֈ��
�7�q�uϟR箘_�C�a�[r+�g�u-'ݯuZg�@��oy�V�5&V�Z�&�(8;��1�2��{k����yo�m�c],Պh4e�)���:�c�,�W�%�� �TZ��tt�f~=$X �ǘxB�ғ�!�U�4������ʫ��:���(xE�#����u����'�x����!Зhy�BI�R�[e�lP��{q H�
��=��n����& ��3B��2ML���� $�іG	��!��[ańāj��o�@�R���h����ɴ�F�;u|@��亻Z�$1������k-�e�nP˧-��]�b���Xbi0xv,nB��2����;�0jn�>e���Ft�.���*f��7\]��,�9�4x�P?:�xf����-׊�j9�8��0���t����U��"?���%k#�P!�Vȍ/[Q3�ɏ�kd�r춂ǳ��� ���ۂ��L�hM4�ʸ���'|�y�0Hj\-{xKvS=���i�]:��a((yW���0�4NMΈ؛�i���밙v'�f��/fH�zΊ�l�'pHW�ً�̑�}Ex����dw���:<_S��\�(���(�����a8���	���]*%/�Ȯ[�����Kb)��$���P�G��� ��Xrw�j�^����Ԛ�]Q��������HRy�$1�$5�{��Q�׹4�Y`��{����G�~�����B򠓘�D/Gj�@n�3~�k�Y{F��d�Scx�\`&\��M��yw���%�h���6���ޖ�!lPi���;:|<�3��ˈ{=�̰�Rk�td��W�'��s�f��B(�y�jc���g�U�3�jV/^�������i�u���kjv?���rAT���0u�cr+	�z� ��6���ˬ&ŬK@���E�l�gDV(g��0LaR�q����yV�SmQ�mH�뼃�=ic�_b(�<��G�4��6W;��u_?� jC�����h �ę-/��2��#Q��f�@0f��x(��j��ms� N�ǚXC�:����D��i�A�:����ݨ�/�b�0Yg��+�]Ʊ���MmO<�|��ߔ]KGҎi//	�f�mjc�85�p���Ȝ����v6���}i1�6Sj�$[�O�-��Z��d��fN3�O�G�
���;����h�^0<�ae����!�z����u�|��K��wr%f�W�C%�[� D�u��z��O� �f); 柃�M$[��Y���V�M����oy�r.����e˻��Qtj�d�g�-��(��d� {�BB�HgJ����`N6O�C��I���]0n@��()bO���1���|G7u�-H�ctn�5{��v���\1�m
���^$���c��9������I�&e��͂U����_����?ĕ��3�m�'(b����΋��:�Q�[ND����z�59r�U��	q�;�іxwۖ�&k($���_v�𛇥Ү:�����\�������7�X��_���Y!0>�fM�G���pn��@4j���&S�=�_!����VX�Me�nrE�Yj"83m��r�#D]��\S�aa�1������uB[ʻQd���i�NP@�p�^�eǎ��N�Ӄ�{��n���ɼ�lY�Խ%�$"a~���b�Y�|�Zci��}�M��Zx��a��Y�׿gq��X��#u����ς��U�ph�|�����L��z�~�Uʪ*E3��y��ݵ7d{��f�Ä���;z/#	-#?[{����N��y*�Ɩܾ��MC� �cA������X��,�U����MB���'�,s� ����v���U/��d4К% ��O%8ԸM:��7+zeA@�4�_Bʯ�z®P�J�/S8�z��h��B�;j������B�!|�Tž����0.�V}6���	R%U!&+Ob:�W������=���ן�ȴ/�����H�f�#��E