XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���eE�����ۚ�*����a.���HB���'��>e�0Q=a��P����ձ��3�C�V@��a����)]� ���=A��a���̰)���9���o�G��=s��'W��s� ��O��E�-h�}:�n�^� ��8�@������i�*�~�FH���ڤ��J��ڀf�%��<%��? T}��Rﬃ���T��:\�ʂ����ed��I&:̉P�������K4�zUH�ZK����t�aC���j���;�0�5��I�y��ɕ�²/q����g����Mh�>���}IOD=�-���m9�a�F�ʉ;�ph-�g����!H�e����fy#�E�7z�'�B��4�R��t�_���݀��/���
�v�	��C��D6��f"yϚ�ĭl:��b.��*�ʅL5��^Sw��<dgkN����{�;W�,|j�����(P9�}*�V��RM�c����7=�BT���qo���[��~�҂��󏕧b��� rIV��0�<k�Eʛ��G��UF���?���Z�V�3���&�	���0��vj� #���a�˞2��!�,�����.KY��\���ta�#�(t���1 .�*���.�5w���9!�]p#	�5��/MW��!���A�#�T����f�њ�~��b.���,ׇ�E?9}�����ʤ����Q����8�
*ʓ�^�b{��a��K�b�!�/,/��@���Ş'XlxVHYEB    fa00    1d70�*q��Uq#e��" E��KL���t�|�Uz.���pvB�Sj�	c	]��u�s,�Z���B�_�!'�ig�)3e@z ��I�J
Y��k����냃'z�5Ieᰯ�\��rOE	�0�-V3���N���C�9�-δ����d�,�E��m��Eh��~��^�?q�_	���'���$z@�)\��_�/��%��R�޷��"֬iBK�t��}��ƃ#�
�{��#����1p�֛DLKw�2�L�oA��^w_P2e���&͔[��?�H��>��>i�R!P'@c���7�DbP2����*�೛Pt*�W_�؍/�����b"��d��o�'2�Ⱥ�M�	�ϩ�������s�i�I_������͑猄��ZȤ`��Ӂ����d+N@�H����E�IOW��Η9�k�W!����g%�a����^�Li�ڛ���ws��<!$G���t�U��#�����6;�z��	��b���PY1}ߜ�S:}Q��O/�|�����J�:�te۔]V#�?V�8$�C�L{ͫw���u�/΂F��w��Kd<h}L���Ui_�4~�<>0�z:Mg�(x��e/B(#��T�y�D#� ]��v���)������*��;*��,����Ԍ@01����M���r/٫�J��W�E�����|�Lg{�GaK��H���<S�`*D��&TC[��oX[�Q�ܞp��>ꉠ�����2��=�D�r�F-�'?J��:s�N�:���wҎ+��Cᬼ��A��g�����1��1��1�@�y\#��;z�E�~-�â��*���~��T.T����?��i,4c�\Ѱ���!̀�w��*CO�*)�ߝ7���T�o�N?��u�ݟ����)}<�%��N��*��8] +:����}�U�t��	��+<#�{v��7	y���x	�8xb����yT� �]:�R�p<��~������`8��2�ڼ����d`�eH��^$�"!@� D�g9�pm���?�61����):qԠ/'k�>H��U5����5��8.<ʹhW�H�)N��ӂe�K��G�+\h"��r���S"�&v{�����D``��ϱI����A	A���~������Tm�E4_���������J_�2fd-���)�l�+s�{�FˑH�?�I��j,#4�lNP���UȦB�F�����)U������mM	�k
����T�����a!�*i�b\-�E2/6��!Uc��C�����G`nu���P7s��D`��(̖��(��-)�$���C�{O�8r!�=�Qj=͑��\�pX����f6��R�-��S�ܔn�5I��Xr��ZF������o�T�m��͈*kh�!�:G�6'J"m��C��ϧ�ys=�x���&4��n%�) )&�:J!�"�ZO��v�a��_�|�'Ӓ����y�`=��?���dT����&Q2�m��B2%�	�@����P��D�`�*	�q@&���W�ӏ
�'F�4v�ʗ�v�FB*<���gE��)o`x��}M��6����BZ��D��Rn��Ƴ �&%@���V��?[KXw�sf�B���;0'ҏ蹞4����b;������X�5�>2�##��'�e��"p[e�Y�O����!���!�|*�#��m�P\���և���T�ڼ������1�H�Ȁ$Ǖ��_~��"�A�򔵎ھS�l��x���
�O��R
�:^d�����8�k<��rBF����b=a��/��O0���p���B�wI��2��>�W�31���:P��C��(^�D�Õ�������.ރ�ā6�UbP�o>L����8��Y]h�Ր�+�r��:�ٜ�=��C�`+�ef׎�w����MQ����;��M�0�X�}�Q^������-6p�w���X��PԚr�x%,�mB��l��?�nc�-H)�&�I~��8\�.�#�&>��CW�D&����M�|X�g�KB��Ȇ�X���D��;��
��R��l������9R�u��Rcp��>�i��)�s�/b�����$��x0#y��a�9��N}������Y�~�*֖&��g��¬V��<�} ^~��h�� 
�b�յ�����9��%��˒Ct�?�!��L�����+�Jw��h��%�#���L��*���/y]�_mD#s<����4i�gP	�~&�xDϹ������k0"c5�S����iU�E���Ƨb��E%���E��v!�s���adBn��^VI���J_ �#E�����Hw���-oI�`�+up?p������7�������P�P��ܶ��N�i���6�ܒ�V��o�{�~�8+���r�Կ8��i�IR��`-aK,�h�+
�M:�׾�r�b70����n���j��T?I� =qɍb�cv�J;iY�T�����#}�v��d=���Pǝ2�2jL�Y(勣��n}�.��GU�ِSɯQEk1���#Z���-��q�$�VἾ2"��B`@��ɹeo�\T��M��
i��EIk--����N-�cEBc�
(�a�e�s'�Coj�3�<^��J�����'��(ri�3��U�r1z)��j�lM!,��Gh!��C)W�τd�N�R�6�Q?xΎ��b���O�5��,I:��H���J��OL��GPV��[��GD	�0�S�����'=����tL���K®�<[��]�����X_�&�m�O�Z�����]��G89��ǽ'���E2�O}r�WKb��nX�<��:�-�Pq���B�����~)�dr��Nh�=~,:����mm�pp�(��H4ߋ� ���,�5�<�>�oȥH`9���:��z���f�~A��&��δ�gŉ'�SG�]��_}��ʷgƒҲ���&Ńuҟ�'2<~����Nɜ�r7���竆��7���)T�s�����I��R���.��۶�]��L�I���v7���Φя��0~�hQ!e��/䗮�9>�~MO�2p�΃��1k�ޟA��|�\���o���@���_Ye&�ac�U�x�D��Ƀ�(�QSݰ��<���%#������RG�����?i#�F�ƒmg<=%��:�~���\/����H*E֒�����<�����W�X�(>���_)�ٔ�!�&3/ �1���]@�(��l>)U�!r�bj���D���;B�LO���1r9u�0���m^�=����ubIG����J:pl���o�>��A-�H����:�T��Q���C)C�l!8���ݡ��刐�i͖���Wa����p$� Cv�1eb��s�h�[J��IE�
��Q�/b֓�g,i�h)���\(Z@-��ǘb=�����bQ�Rۅ�t'�?��ۮ7Z�vx�En ��i��o�$�aJ	b)lqY�F|������te�a��I�%���_��Y+���A)�?6%mȚ�W��ֹdA��_��$">��ެ<3ʍS�`:Cv
���j��_4�J�T�)�������/L�x�Y���M�k,�z<��+� �vl��9?C^ts>��A�[uXO��oęǆ�]�/Tal���s� �������?��]��a��&����#����i2F����%+�����v&�מ�?�8���	P]��<��c����`AV�Ys5��3�V��AJ����Zw����i�]�ZPhI4���JW���5�&Ԁ���V�\_mgr\��an2O�&4�.*5�DY�PKѴ�9��cX����7�2}�|j�H�	��̚�);�|+��D���j�'��N7�{U?��n��b����2U�I��bc��ĩZ��J�8Y��,im]3�o�H��K���	�lC>�G����E�Jhg}<�Z</N�Q����Q�&� @��S`�j�O��/X�r�S���N, T7MŎ��cK���UgN�X��Q�L�t$[!�+(t}<p�ǘ�4�;ȉ�۱�W�
��h��xk
X�Y�Z���G��KN*���'ҩ}�w�3D(�3����a�ǛU{�sy�[��eI��B]��WKV��'��
]�;�X�v��)�����3��~d�zT)�@p|�>��$R�cy�¾6�ɌL��h茦3}!0�6�[�������U�^�:'��͍b�v �Y}�d����Z��nO�S�Lr�������}�ʨe'`���h�Uq���������c:�PB.~���Ta}͞�*��n���;�|��/���(a�m��Ҝ�3	�q+e�f�P��r�#�e�*ގ탦��\֕$�;�d�p�̸�� ioZJ���;����F_�i��ɭ\.B�
s��b
:��q���z5��f#&Y��Zx���y�j��J���#1��·l���3�r����Q)�E�h�v��R0e:3J]0P@��J�0������� �����wFs0v�dsږ���U�����q����I���SF���)��O��8<�v�z��Q5(zO)��"9?��U�N��@\e�>/�R(���gR2��	���9�S��}l����,T�7bM#fq��j�]�9��+�9��g�ܜ�y�5dc�,O��f�[,�M�;���F�ↄ�Y�*5P�˂&F�'��Ue�&�[�j���"g�݆ �����2���v��WdM����!��/��e�_��Q��+�ޯ�a���dy7FBD�RC�����/��0!��\pp�E,����c��^���!m��n�7��A�*ԌbA-9.��=U��J!�,���I�G��ǋ�lܔ�C�&��g�:��3}�4qM��oM�d�O��): ���������C���dʶ"�S��0 0�j�N�m�S��?�yY'R������!ÞІ�/��W�5!���~�~� Mg~�������z@F��]�$� !�?�I����u� �#�f�H�j9�h��?W�7��P��<�wsnmz���2���6-p�b�@`{J�)�eX��A6˄��b.�M��/U����,4����=N��^H��y^������2c�o�Z�Bۼ��-���2~1�ϽW��.����>)��)geaK���Q�&����=eiF��:��nG��V��3/�2I�be�l$}) �:���T����angm1�L��z�GB+r(��yE�j�&R=ۖ�D!��lB�e� iv�<K]|�ty�������)9��ܓ���
��n�0�j�W����a1��n>޼��7��2�e�� �����Fn��C)�D^U��e[�H�<��?)�*�+טk.T>\?r4V�e/b�}n9�a����_XA׶q~�x����[���|�F&m?���޻w�i���tr��߬��1�1+����qd!��>?o$��˵�bA;/��ù�2>c�e���2����5����5%���Υ�����j'H ؕ�^��T�;�oX�Ģ�X�a�⁕ {1�1���!��(Lu��W���7�����:�-wۺ����_��L��X��$���E�`UT���������l��%���|��,g������4��6iu���s�D��_�L�� ($�iA�ވ;X�}?��b���h���v���ߴ�w�
� �`@wm�N��b�I�������T�m�:�~`[���Ţ�v^�A*�.�mѸd���ye�t���jT܆����7�;�1H�����d.�ʨ�P�b�p�����7J��m@U�^h����I�-�����w���j$Ƙs�1��8���ˡxc�<K)��g�}Q�����'5�R˹����>J6%�g9���9�mb��e��Qc;x>���י,�=��A^4�tR	z�}�S� ����!����|R$��N\�!�G���ހ���I�d%r*�T7=��!�8�A�
�8.�@���X�'�"��,`�=uh_�gE�/̟{7�e]�#�a:D��DN��K�1�(�]��,��N���`J�9��	Q���5����l	���\0pė~ �b ����*�T>�mY}�#U�� `B��M�C�������Z+��������Eϫ�y�񑒜z�H쳕���τ�`}�^��P�(�}O��L3�y�c��Y��$��(����ӊ������Ζ�A���Z温���0;�[!�ˈD��zL�η�bz�[lR�s�����`���um��YX�f"1VI��_lW�~F�֋'�&%e�i:+�o�����y���j�T�pY-[Vh��h�D��]�h_[�]�����l^�A���}n�F�O�LѾJ�yV?�1�GB����$�{�Lm<�t�.+mHʍR?�q��`�d���}}�]q]�q�Ʋ�I�J,J7�ɎklF��`.uD�z�a~��U�t��פ��Gɶ�/K�V2!\�c�j>۽�#�KG���16����$�c��Z)�70��-�^z�i	�r�m=�?T�`�	��CO�m��
���^UM3��<T���/�ޗÊ��@KMjN��z��
�/��w� ��T	E�(��Rڂ�N�����l0��h6�R��mf5�;���W����B9�}
mq�cJ�"q��B�P�sH�=Tp���!8,����a���pyj���MR�j\��4��ɺ/QR;�,*�A���+��j��Dtؑ�|��1㬶��LE�5s[2�P�曩"[��M�sѺo�MT��AHĻ�k��px��~��3����_EG������=C�_��`�������2��]���]T"JF5�Fg��]��/�5�@DR[�&�WQ^��������S�?"�^�cypq���w�Zbr��KK-�>܋Uq��(*�=S����_�C���Վ�(�c������=\_널��0��u�ٯ��\ߖ��@h�;{_��r�N�W���T��(�g���b� �(�9�	L��p�����6d�k {:6�������Q���l.,ԓ8}��0��s2'�
u돠��0��B۔_߼��:rr��?q,J����p�-�þ	�o�,C�߸�$n����&ŽdE�����hؘ�6��a�;!��0�8c�z@��<���[�9$By<� 8$�vV\�)�� ��<�_cy�9ɋĶ��C�6��V}�SOa�� 0��#��Zl(��W�z"�n��ר8@M
u�f%m%ڱ�<�''m���7�x�����qL�+3��BXv��4�<=茅���@Oi� �x0p!/}����<�O��"$2-�՟Q�� �OIȗq�B�z���Hs��L�Vd��୦�R��/�;9�Zr 3�Шm�X��©��vo��\�p����u�r����Ҭ޷|���,DU���������6��F"�۷�Y+��24?{��aTi��Ň�˄I��B@�l/��ň�v�Q7#^ffb�|U�.�8�=ͺ����cC��K�cKv�?r��XlxVHYEB    22d3     6b0��.��҇��٥U������o��8�tDt�-�7��S�4�&���Y�.��FDXhӉ�j%g�V���}�gޡT�������1Ƣ��9�I��f�s��DV��M�1T���l�n�}&@}�|@�?��`�@�3�zicԺY��5/�x���%���,�-½�C�!M�D�%J��3.��a�����8��u� .����4�M��8�:������|[���,!8�aX���Qqw�E���Mb�I'}�}%��}jE%�v~^S�Ij��o%;����&܍@���b����P��K3C�x���S�43��N��|[����`P�w ѽ,iQxb"�&Ҝ]���s�D���O������$y�A燥>N�jP-��YK)��x�y��!�Wt�{C��"�v *+�̅�KJZP7��*�
���f0�ș����av\��@�`�,w�����9tN�A���N����e9��^XO���Ŀ�+%�;�v��(e��eE1�'%pn}�*���8�n&LBL	���,�����ŏ@��ݴq×����Z�:�K��G�j>�Ͻ@����w��3��H�F=�i���x����L kd@*�0_?��3!��'ev1��wÙ�bh�=Ej�e�*�P
o�{_q4��U�D�Z3 EPS��k4'IqpH����ZP��R�����Ö.�x����*�lk����K�㓿d�E����d%��2��9����z��¶�C��s�C�%�@�<�HP)	i�'�������.�OӮ!k;���y�P�5]�VMT�/�]�2[-'v3J�{3�������7��;O\�ee�=�w�H�]��h����.S)���O7tG�{+��/�����[�#5�|ͼ�|6ǖ��J/Tf�2in���oti@8�Y'�[���^��F���
X�,��MEh��آ��?�B%�*Ş7B�)�����`?��%�'FֶnnfCf�- AY� <���R��c�z^��=Y�����ja�j��� *W��\C��s�>��gr�y�rџ��L�{1n���Q��~�1���>S�ӟM��<�2�R_O^�Ju���|?9[:�l<QS���iv�ǌ��P�h�-���1�C��U.s`�]�+�P������0+��J�͗�b�C}@.�lF�Rz��U�tk�h���q�ҡj�&����a�	J���t�\GFUT�O{��ƙE
��6���JOtq�]w[�2�d�L����_���P+�s�����oЀ��p&�q�X�.}T�-?���7*�=�W���)r�~s~�x�ў����$BR2<ڋ%��d�H@�\�����U�=�$�2�S��4����q8
�c*OʜF��kP�*��m�"2�;������>�{�*w#�d:�.�g��ص:�(A)�r�ď��0"8����V��F,փ��W�uRkSJ</���XmS��;[�_l����8U����`���X�I��,���d?/�G;.{a�R�ۋ�4�֤l=�����9fٷi��*�d<�������ɚ��o"��v���f���C^�7|�o��OwXI�ˈV�o���5�ۻ��Kz.\'d� ?�v(�C�eP!�"��o����[�/(�����dB�r��=�ֹ`���Wt�U��e�����A�kW.