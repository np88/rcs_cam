XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��F|e�>m	հaC	Pt	�
��`�v\6��Kc�K�g��)?����$yi��E�.�-r�j8�y��L��S���� �q�d	��e,���Z��U����7�X~��������y/�w��o���]�cY��Ɋxq$( ��D�-� �H1qf�a�#���.eݍ���39��/q��l[,W�J�%:���&b�F�P��~�T)��)�.���ڍ|S��:pJ�񿕵gQ��wJ,V��o[lYm/-8���;,�!�fL���s,ӕ�%)��2q�{6y�$n���*>���}�� ̘�-}I�<T�wf�������t:y�C��^��^�L���Lj� 0y9����d
gX��"!q���v9�DY]u�Q��m�VH�I�O���;�M`b�YX�|GE��i��۩�m*ɣ�ʂ[A�t�a��y��!�*A˅�yI����Ж�w�j��*!�_Ya���S��?I��RG2#�LH����_�V�T~N��H�C���O�<��;�c^���؋�~w<*t� A�p��~���-�h!��4�@� ��*Q�k��\{oC�ܹz��mъ�Sڀ�n���gc���?�2�2�JѮ��A�=�HX���X�P��<v�0(�򀛸}�4����%.�u;)���&Kr�6~D(���#+�UZ3ŷҰ �&�~�0/����l�Ov
D~��/��\��VaZ��g*Fc��s�V��a��H c���JQ F�+,Fb�L�7��XlxVHYEB    7744    1780U�ڕ..�����U�ɶ�� ���@������в��W�E�Ln�MB
���&[+�h�B(�c����lW[��c����W\`c�j�DD�Z�n�1��ۀ�dGÈ�%�޹
?��S��9�^a9����E�Cy�|��&F�`��j뽪*��w�bc��c��)�s�UvJ�v�3`\4�
��;������G��O����!c}�.��w�u31"&�Y�71%:������~L��G���ԇ�7d��K	*ĽH�h4�����_u�JD*��8�:�vY��W	D������<��Lw�.I%f%{ ��v6�,�Jl`Z�ؾ^�3͑�_��ֻF����e� �H񅉥���� 	7	�m���\���V���=��A���N�t�G���VY47�I7/�F�I� ���	���I �Mb%�4aa;j#�F�<8�8^�Y,�]ZN�C��/�(|�F�A�&�Sz�I�(zߓn�9Q��m�����"%���lIIUV,�3*��ɦ��@�7D4�sb�����6	�|XD2b��q�rs�_%�5��Jɟ�fV��Hu�y���amWo� b����?
��|U@�"�`�������L�F��'�H����VD����������km���O{`�� ���F�͠�4&�Q(5f�s&���fUW��ԗ\5�/R��WT�Z
S/Ͳ(b(�j;\&n�KH~LD��P���5������'���J]z�
C��K%�mz{}J���!2#S��~��YWݏ�K��w���d2\G#��C�F^�;�r��������L���Њ��P��2��0�@���i-e��o�(a�U�c'��J�N?Q�mз���@�eZ}^�L�p�Bvѿ����#p��L}�ۏ>��i�Cq��K�"���r���%���ͦ���0��ʜ>�iM帏�H����B7�<�mma@l�o�#u,�`��V�?�;9�������\ˇQ���W8ʝ����K1X���*�kx>$��У�	���_N�v�a�/u����s�.���ד��L�U��v��Y���4�Qa�H�>8���M�`^����("�`iB�L��	[>���_J�Kv��ef���B�����[wɌ�xB-z��xaa-XmZ�K9�<u1��m(9����0��~�������a��1�"��g딈���w"�X����#�#���*�~��yIA�u�ㅨ+�o`.l[.�xzY'�s)i4�ee��%�~���pmh��D��w��3�p���nP��N�u�<Q;{��'d���. .ȿ���/�,�yV;X4f��!��E�6fD�{���v���N�*$�����@Mx_�C�*�0}ytqW���Ovbvo�b�(&�W��c�c}���{�-��5ӏ��8a���&G�h�A�	�GV��ġ�q�Y���ۏT���c�r� �����+̴��=��5�M�f��;WR�ˠ�K�Tg�i���+&�n���5��ΓoZ)<|�u��']���X+߷��=v��k����g�Pk�q��52�`��S0`�-���t�жy6��	�y����l�F'��Щ� ��J�k�"e��;j�Z�����_�̍�FU�t1S��I�FD3�9>i��`յ��0�r2����G�f_t���M�oM�5�J�98��V�" ���r�Q�&�n2\~��z�.P)Ǌ!��@��>|FFF�ǀ��M�F��N�*)��+�[0����3FC[,�!��t�Ehɕ��`���<;��S�5�p�@�����]"8J3��󻂿�}w�ߗ[(�?��}�G�*��y��ά�8�r�_�9��4���bt���%ORq(܂���<3#V��T�h��ߔ�*X:�K|�7�{�E�+ܠ=ME"���0E/��r��Ws�8^+�q?���B*��X=P�MND��Z�YqE��_id�����E��C�9��u�+&��� �5�}�/���!��+�h��h<�	Ӧj�ÕڸTN'�5�M�U4�
/�n��x!M�2��G�@�D���Jq�_/$�QN^Ύ[���MG�~��.��*�"oo��	D�%6�:�.���C=���܍��U����z��O���W�೛'�p�#W��ϋ��|]W�X-iͮ�R{Q��.�a6���'�.�Y:�)Kq�,��Z�I��>;��9��[�(�R.��;�c}�J�"�-Z�,i�ϙLG[R����ز�I��)�xM?q���1j���vɮ�ϾBX���A�w�n��� H�6��:�J�����@E٢���h_$�"x��0e(���@XB��F�@��^~�MB�D�qw�ċ9+"��\���^ol�]=on��Ү��p2]�]z��r������j��r�+d�����$�m�Ni�Px!&e���]��I�k�D�� ��["���H}�4��,5MX���HHV�{�㫌�bY?�h���}cq��3�?� �g�bVA{4��C&Ϊ���.:�p�qb�:�&|�6�\tϱ����/�*i��=�KG��|���ՉI��N�y�!�]cQ�_6u����R�0�
�u���r��z㍝��J�e��D��B���L�Fݗֲ�gӜcH�T�R��r�Ϳ�晔�/a����0�.2����1��g����٭o����!	VuV�����ŵ�fm����2�I<]d2qeY�"�*��\T{���L����UL�Dǐ�N�ILU�nR��}��ky^)&K-�+�n�#?((����rdXǽl�l��~�����R�����'k�R��1g�K��gڬ+��K^Q��Xћ�mQ�f��H��@	��S]]��ȍ�4�T�y_�#y��jP���@���A(��ԗ���b{n��a^%o�\ϑR�Yŭ2��c9�� aEm�Z���4G�&�MbFz��UF�A�X&��-Պ^���X�����@�tt�M�XgX�nE~Ʌ1� �X)�b��rM�L�
3,���Zv5�7���NrP�F�wxS���Q��0���L\#/
y�2����6�-��g9�*��r6gqd��`�^]��N��U�舍˚� �I`�ɐf�3Rh2�ňN�o���a�xQUr��D#�c�cTS,�1��\�fM������g"�ekuLP	B�&s��a��{�(������\�z�1^	�/:�"H���&�z�tb�<��"�tf�=izC����2JDE�#~r���=�~���Q\��G�x�>W0k?��:�rP�`5�@��A�/����+�X�(b-? qg��"��dwwE���Z~�^x�Gk����W�����8-c��@�ٴi����19���4���\��$�����dg��uMڪ0	���Z�R3?�"S<�_d���5�$M�o�q�`ۛ����c�`�]6��څ�@�Lٗ���aj�P���d�kE�b�DK�Ezk_�A
��x���q�2f
d�r�^Su<�|����׻�hw�a��G��'eZ<|���h�Tw��LH�/��4Ռ%�#�<Gl�.�A�S�8���K��'9��+W�����L���ˡ����S_�2��;}��-�ת�sC�]�S`��0�� ��Ͽ��Eﬦ����k��w��!���U�;
^�_Hɺ�f��"R�+#��|����~��"�a�t;��(���c��%�������E݌�%l��-lO�co���x�[�	�O�O
4΃�;��|N��G���t��?j.���%�HŽ�A��QW���D[I-#�{�׺���K�P�,���"ƪ��JhòY�z���õ��s��a��w��2��|�|Bp�p��e4��f�Wk�F@A����[G��GL�u5�iW!'�53����L�#m#+�ܚԌ�ܩ!��tP\P�E��t�`�L�7���:D�SP}�!0��!
I��KQhM�3ԧ�gf>0�E-�����=T�n߲�võ��:eL����Ξ"��\��j��v��63U�����h�}m��h|*�5��zsYD����_��&/�c�q��u��yJ����LqǑ�Cá�A�Jh�o���AH>���STc7A�bL���xZ/I��W@W���^�����ŚhFI6�f�$n-��~�'V�
��Ro#��$�l��LHo��.Ρ�̸E���.?�t��;��S��e�ĉ ]�x��__>�3���)���¡:��U��r�N;\�[G	,�x��S8]ȍ�{T�M-��������j�_��'��|���크H�-o%������ANh�ֵsˌ��7�]�du���z�#U�}&���?�l�cR[#F�HR��pub�U�����K�p4��J�V����Vz�[,��v����<��#�8f�lزu��i,F��F�f3��7?�G�L/w�DWGT$�\n3��B�V��Nx8`?p�3]QJ��b�7�-��nVxxDW�9��R>{@�s�3;���
S�n>�f�:�)�r��몆״U��WأfW�<م!S��Y������W����#��፶S�m�7t�{��w����Xlu�#��B�۾����3�a?���?��"�s���~w��;|���7��d"-��� ��M��8[k���A�$�֡3';�N4�����@t�1.a���)l���X����$	
��V�3�A�=A�9���i����3G�����%3[̎��Ss�7T�v\͌�z=���_�}����F7Pc��s7��Z�YR�?C�x��@(U�;[NgH���װ��Ȟ���'�͡�$cf� P�y�;��V&9\xp�<� � �4�AK:�a{ l)
P��/�~/&� �f5��h&Z)�yu�O�8e�E���dQ��؁b�{ǋ�5� ��Ȥ:G�*Ń���n{��	��^skN��.�h��<���at��7j�P:՛�@{������`/Q�|zj:=�I������w*(�@����Xu��7'�\�(�P��7�Xk�/7ˌ�F�-�6�H�_��~�P�{���O�<IX��N�{9
���o�0��;���j۫�q5����Ze6{�v	O.�>��Xo�� ��%Z-���+��B�8d��@�-�W�i����6�,(���N̠��@L�FO!�_�*�r��6����]����%d�P&�+�������QT�ꅁ�̘�a�=�pη�o�
}�-���L�fwѕQ�d��J�H���&���ԐU~�	�dҴ#WO�";en\�#����?�?��<X{��h����毀��0(
�Wo�Qݸ���)�k�wL��,��oXI���,��ډ�Ż�ZG�fa�V�qRs�+��#X��l���u����z�(�p6�8B�H�G�����
V]�`zz����X �y��R���*��l��P7'q�1���]a��>{���$�Q��AAr7�Q�G��$��B��g!����Ԫ$�7���!��yb}]�|�.�}?�m젺���e%�Ųڲ]+��*r�;�HE%ʧ���9x~JM��1��|[6F�%�$�	�����ZA��K��KpH���/M��d�z���ŧ���["�O�;�%��Ѭ�3ܐ�:	' }���>��Ԑ���"�}�ڎƗ��)wy�@B��}8�Ї�/Ô���i��t[؀	|̈́�LHV^StX��1�qK�v�y�*�Qzj훥��~Ǆ/l�Az���8�����W�튬��!*�T�冾;Μ25�g��^�WhzFF3��pP�6?0�&=;1z�/�z�A��JѾIq��(2]0;�2u�Yzn(����u�����=�@�bk����/�,�Q�����M�" ���5�UxѰ.D�ܸ�����w��Y͵�I�:|���]�k�$�ap�|t��������7��,�m(FA� =���iͤ���l�d���L|��|�Ƀ�Ԁ�WW%��D��!U\�