XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����3?!�t���4:]�y��A��'�ϼ���=����8�{|���50�m�6D��.F�g$�5��>��TS*��T���t�D��/'�mz*�����ݠ@3�6�g{��p��\Ɩ�Y�c���$�\��R���ϥ�+.�Z�������X+��;.�����d`)틢r�<"&�	Z����CA�J;&D	
��*��bB�L�5�H�ן�bh Ԭ'��+�;���N�@B���U�l,m~c�-A�&O�����@*c�3L�����{L,�y�U��rN�QTcXVË�5�)y]�,s�'��>¢Jzx���U�5@t�7nI}�끊C�&zۊ�6�y?������n�a�m�A6@G�	�⏙��zþƀ����A���42��Ѡ�;�PN=9���b.�B%��^W5�X.��:�Y�	qE\�d/(N������̃Ș�,$�C�&�^������'ci�d�����<K�1C�XF��( �	��DVK���<� 52Tv=�.���ޡ�U��R��`7�8\Ĩ!�<��g�:f���j�Eb���ӆ<���>6���6�י�����f�n;���g���0�ٔ���>f�V>���me�j7����ͼ��N��2����Ħ�P�%�I��aݮ���4}�
w*�~
�L��9{�j�RQ���>f(�����#�F�+���{�O`7A�'�)3�ɼ��B)�b������3��T2�H�e�d	��'i.E�6XlxVHYEB    3099     c40�ƚm]���>��WQ2�܍�����s��b���P�K4�i�OY#xR61���$��B���Jԍq�Lh�Kf+�:��wU�w��!:<���I0o(i,֘��0���s��Y]w�Ƀ;��bb�|����!��l���8��0vC�t_J�4���2�T�5g�i�\(�iV����v�ro�H�!��"�~�c�.�
HP�V���Q�w�r^�$j��)���<�>8�X|Hb��P��G�~3y�p�Z+�ա��`˰�E����j�� Үݳ�]`M���>Mx1���!��t�Lj|�h�4a%�ɬ�s;�	���[�,��>��,ln��`��g���C �<�o��ٖ_���XƿUJxb���5q��Zu+@ky��J��x
�C5P�p�E6����Wm(	%�\!�d8a���
)Z#A��P6XA��%-��1�.�S:���
iӝiM�1_��9��g����9�pEÄQ�RM|����r��o�y�lM�fp̷�X�5g��v�:�c�#��@A�@���-�Lf&�aU��^��cbx�'�h��*��,3�\���IIX×�L��!��O��'���VP�e�� ��,zH3� H!5e�u�3�h�Z4NU.cC� ~���|B�AX�k!��t�R@я�в���! ;�F׃���8"��zޓi.o��U��Ib�X�Ƚ	�R^�����Õ��|�Y�U+[֢��@�zKv��	��I��V�nN���<��ΰ�ۮ��o�L�D�{��Ҡ�ÉLS:0b,@N���mΐ:"Z��V�w"y�q�k^���UMVf��a�.�p��%}�&8 %�e)�бSwT�-�릴�1o���Ǐ/���i����}�va�N��#��.r���$��Bn1�&�B �xET�=�իx�Y�:���>��\��5�lK�@�/�Lw�XR 
#����ј��4��y7�I��e���9G���U)0�L:��x���z&����-���]��X���B�����+^�^U�ګG��u� F>�#�	�w�cMaa%�u�����=D���=P9ߺ|�x7�����\	Ci���r��Ix�d'fخ(>���5�6���9y?n��I��(��d'��Dǘ����)pB���cJH���7ع�Y���1����&P\;d����a����������3M�z�r'�����&	�%�c� �I;&��]�m�A�6��Y3�o6����<%t�.�5K�	vJ~��|��w߄iŢ��o�~�a���bP������.��GN��:�F��Ҍbx����1�&M���C&��7vB�Y�<�գ�-]Z�'%��qEE4��e����S�O���֬BՍ���W�3��/9(Ae�kw��@���J��<��Ղ����&��1�F�,�G�}&��=�O��a}��D��H�bM�ɤ?�{���:�U`1���̊����F�܇9�o}AF� ������O�*�M��Q
�#���W)kZX���@%�%-��q�ﵩbgLwP&��=�x2ߕ_��Up��@>_&�!+�����\���n���  Kq-9��l�;�E���0`:��RՀL��U�Y)�)ֳ��p�kP�cp�(*y�,R$�8 JXD�^#K(t��9�֭XCX�
�Q����}�?�����%X� ��j*�����k��#̆��6����)~�귲��c|�����.*9��=�j=�-'�ɸ�B�5�B�/nWI�&�&�I\��o�՟�:����ˈ��:D����u�Ip	���6��02����R��\��7C$��#>���D74�A��ܹ�.}sđ�������+����_�%l�fv��CKd&D���\(x�.��O����[]���W�p6��Ng׸2��]H��QR�%�j�-��@�^��I�@C8;/�{�yZWX���a��q�1�s{A$��&8Ž�j 3֫���m��@�t�ꐖ?�c�Di�Ĭ*��u�	u��{���3j�/
<���:=�O����9��۸}�9��t���;�RL�?볯��!����7�`zǜ�_�\^] �}����*��Y[�\������v*�fO�U��[���]�4���gr�����R�|���ne/�
�hcO;h� �W�����A�%RL��R�Q���V����i�YsU	0���X�qb��u�,+�9�k���]W�&t�yU<m��Ax�*̒�+'{�ۿ�W��j���I��`�yL�)K�sk_5��0����	s��C����l�A,����y�Y�[�Ð���Z	78�-952�+��9d���
^զm
���J ?NS2ܿyu
%��%�n�䍾8�k^�&Ǥ��Y�I���=h���VLq>(i�T�p�4��0�e��!	5���S/5���r[9g���	I_G�� ��@i�P.�DO�ڝ�NOg\)^r�u�Vb���ȑ�H^q��S��8/n�=3��揽�{$��ɹ���候�B���� Ǔ��:��'l�"+���,>y��t�� %2���°������\e�G�-Sj٭:�)~� ���-�:7YeЋP�v� ��B����L'�E������!y���[C�=���"2��.|����O��9��5?Z(��K,�"S�xYW�����V�K�a��x�1�Kr21;��~,��ۏ���~27΂g�?��5Ӎ�09�"�A,6��Ķ���W�)Ǳl�|���/RCr��Q.��_k��Xʥ�;�q���<��?j�^�s�-��]c�\z=�o����L]M��4F�	��8*���r:,����7�;������i�K�PI��S�����o`����j�:��\� ��������ۡ�^4N`�j�Д�vHߞ�b��F^ҷ�ٯ�C���4���Y�Jo|x�m|�x;{��`���H��Þ ����|���h���C:E=�XL?�4�E�R�;�j�3r]O�Hl�(.	vPj�XTE����[X�=M�~&G��
jo�ȩ.L!O��!g���1A��t�b����c-Z
@5R��H>����a���3qU,�\U��$��[pV��L±��;�5�k�WA����7���