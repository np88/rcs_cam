XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����C�(ē]�5=��j������H'�ݴ�/,��E��=|mLa3�s1��}�Q>j�1b<�����cҟ� ��U2Js�̩�$o��>r4j.����|R���f�O�]KQK�-O�U�N&���f㠱���A'E�c�>��=.F��<_��=��yf&�t��!^��-�k2��zș�z�X�r�i�jq̬�O]�SJr �1?#�^�	{Z}�|���M��$�E�3�F�l4����$U���4�u��r)�cZXQ�;�U�,�Ym 	�;{z�W��?�tO8O%��B�N��)��6���H�F�6��PFl�R?��r��sH���I������hu���z�9?TZC#_ BDs�s�5��pB$\3�wĀ�!��x�85�h7�B��pĺ�FL���b�
.;�=�F���Ԯ��Z*:wVU���(?���7�o
������;��1��}ӗ=��O�������꽐4ڛ��%���f���8��6;E���ݙ߯S+S�Z�aY��sw!��9ͻU�*���z�"n��J�p2�K3F9���	�g$�C���@�j�ܐ��]3��:F�#�(	~�4|�Y�������m���US�g�����!5�Ww��E@@Q�HԹ/6k�J�����_P�jT�ec`������c�=��T1UCg���(8y6��7.����\�N��&�GU�Ϳժ�	{��wGv�����������5��2�39�ևf��BeT�9g��XlxVHYEB    162c     850I�}�>�/k_�BC�ڧ4�>K|��г��S�}�K�n
�0`Ss����1G���L5_���F��j�Os6����q������)-�ku߷���U�Qn����;�E=��s�]�hJ�_c�ES����Ѳu�DΙ�3�]}T����ֶ��9���� ֐yÏ(u`R�"4dR�@�����+5�#����沃�o��l,�K��P�&��k�po 4���y� �����Į��2����\2���"qيiA�̡�ٱ��%�0�ܽ;��*�n�-s�n+i&u�x�H��$M�;^	��B�ů�yvn!�f�6����g�� 9��^�Z5a �lhJ�����+S��Y��rb��EW�^o�/п�6��f��U��d[O�'��`�٨� �����C�z!\�=��_�۔T<м����D�dY�%`������*(���]��.#SAe�R����Y>���a �@"�H�>޷�g�.l��*Giq�PJ�&�{�2݂�C�YMB��`Wc�l��%�0�6�M���Ž��a'�d��^ Dya��b� ���j1xa��9��Gl�os}/5�+8&>td<�.D��;uE�L�	UĮ�.ٰd!�ç�״��`��w��X�0�� P���¬�PT���t�~:[��n���/��R�.A�,�kaCNqb���A���a�8 �~����+[�N�dD���p�vh6=�!��3IM���j _V�(B<O�@�:/⩢�]�St�:�JB��~t��Dz�r���H�HJ�O�ݒ4q�.^�$�o���v.r�G��T��3� ;��vEqe�~X����E��^�D���\��ˬ
&�4:���o�X4_����Z��hn�a�ЕR���^��[�a�=�EZ��oi<�^0�W9����n�k����&LrW�{���dg032]�VGֈRD�Y��z��a#��Jl�����{}��ߌ�G@��z�Xn*�&��vB������8�A�U��4��>�,�s��֪�;��^P�܌ ny��v~�*Z��WO�LF�����	eq�W�>�uczoUA#m����Z�t�����e������d\%_ZP���b]�p����do"��
Ri���4A{�y���]�k6H������Is"�ru��-b��Wf�I#��;w�Y]�������jeA�mHso�vp���g��a���S���G?a���:^�4���#��UY/
�ab+��i�ӄ�ߛL�p�Y ��b>�i�?�}�����3P�t���(Qk��G5L�^�M��d��m�>&�5w�����I>��ӹ��:�5���%��
�PX�0q�X��V�46E��rحT������<�V��Z�Z$�k�h��;���<O�v�V�.�@#��SB�'��Jac;Ӟ� ���}�c��� � ��,�3U�N�[������w�X�m{���n���M���Ȼ��.E��D��]hu��g;"�t��9ɺ��~�Q���2�+�u��0d��c
�7��1א�yMCu�ס/��#����|p���:ΟZ)�7~���
�U!U����h�mh3���MZu%qj���tp����	*E�皚ޒ����+�r��%��-���-zh^g��Zr.�p�u�@���V7����Ҙ3H�8ΰ���qB*�u/J�x���$[�#���/�8���,��\�}���\�1���KD��0��1b���e@�t�r7��Vyj�T�0��ah��V�v�x��B]��X_땆��P�Ћ ���O�k�|�m��%I��?Sdd�0�3̼ ���O&�|f�vC�*R���ͷ��u;�ۘʙ�Gœ�M�8`d�@3���
<�f�5;��S ��;ǚ]�a��ks1Q7�R+M�P���:u|W/Qh(zz�u�sP�q��Ñ�	!�����X�ooA�6�J\3r�7�|y���W �T���}�<Uc�4Y����aã����s�2���CV��^�MRr���/)�iSifݖ�� Ӌ��ԭAy}��_:(;f~��	��e%<�d��B��Q����9h�a�-����Ҁ��=����'r+בXH޾�ץ