XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����`�E!�?h�v��e,����G�D�j�^��8��*��@��A�6�o�~[��e����r��{�F������(��
t�ts���l����	!���[�P���2�-#���R�A�-��[��2��/u,��Ŋ�p�}�W���dRP���t�P=G����~���q��{�:�1�D�"u�J&J%����[pɳ�O�Hݻ�'�L:E7\#%:_��SG�z�"|����^��MQd��y��Z��J�:�]&�J���y�k�ѽȆ0��ț�f�B�P�W���|����x���ڿ	�Y�J�A����<)էբgv��56���֧�xT���)UsŤ�	���k���k�ɜ�φ�i�̑��@�UQ�z�����nwa-�Ҁo��Y�}��/�T�%��y� �u���cg	�&��׾�� 6 �óqS-����=���ԅ��cC�x<��v����M'�j�Jy�P����r�ņ�$q���=�;�Px��f�x��Tfy]^���L8�a2u��?un��.W���Z;r��R%���]֮��%8�-�7T9X��6l���=�~���� ��<Lj��� ,�<U+s�t|n=jf ���SI��ejy��*��^����xyi�+צ� �C��NBjf��a+y�fp@)񊄑'J7dT�����د1�3[�sy}3�\�}}9x,0#����ɚe���� s��V���v
j��|pb�7q ��;�{q@�G|d�tcO�w�ّ�����XlxVHYEB    b8a6    1ac0j۹��b6v�5��h��Țx�Q,�_��QH�������)�A��d�f���/!�9��W褞ܖ��k������ـX�prG���-���2����!�щ����ȪT�T�ݧ]�����6��s�XN3�JT����=���}e/o���u��?��d�t�e$S�-�&?����~v��L9 bɲ{3�7b�v�� �q�1��4�@E���+��K6N�9��.�Rn+�
��n����Y{��4���}-��	�iL',t��c���1���V�1Ou�n{if�0�?���<�m?�rT���q����Z򼽌��~h��^d�_�bR�J�9Fk�"�Ӱ��H�`�R��g�H��hE����������$'T���u�W�(��\B.Ns���I����:���S4Jt��iG��Juh���{��n�Zu��Q��hk�ǈ���Tn��E���L�c�8o�|\���F	�Q�~�htx0l����5�پŧ�rgc�>l#�k)���*u�0�ܝ�װ��!P�E��F>��̎{��O��7g�Xo�A�{��:��G�u��6�v���er2К�����DAf$o�"PX�rF�ނy���aYx]�s�v84��QT�O	tC����C+��Z���a�;c�bO1�u������b�,M�9�ujV�� 7�jDr��s���kk)?��'y�v�!*e%�����>/d�5���X�;��kUj~Hݷ�j��Q	��$�AU=��HhO���G|C>�K/�g��4e�!�D�o'�1؇�v�cЌN�q߂��td�*�5ٽ9�W��?��������D����L�M�\��5��.��G����E�Y`�9�=k�h��	R�j�<���=D)i|8nH�b�Lf�ɩ��0�O���rK���N�����oN�;��2�>D�D�Rz�:�i�ʗ�	�|�؎�P�U��k9�TY�$�H߆�ra� �.�u�A@y�a�G�m�<�����R�\y׮R?8��c"P�>�\z��~BX���)?Գ����A�t�Z�����x��?��"#4��6�8y�����-m�)i�Ѻˍ0\� ���jo{���tWg#��zE�J`p������E�<H�c�Au��ʦ4����s	���c{K/�u�z�
4p\���olS�m)���81ى�y7�}��5�9�"�̓iҹ�~���n/l�4n�A�Xi���1�5��Ɠ��Ul�����`��4}�{�S�W���i�|����ep�x�=�b��b	��%6Ğ�=�^}X[3-�s��#1=�)_c��l�65tM<�R���S��vŕ���^�^'}m#,�64[�}ԅ5Y2���Z��/aUi����G!H��zpP��)hu��4�,f���$G(�Θi^��8�U�����!�eD��BߍoB�o<Ao�#��N!�	Q#����vT�f�?[)�.��(�8����o��E��җ;�k:���W�(�7�$��f�;|r�R`씉����<�d��d��绣k�wtTgC}�����'j��������pT�s~�n��f˥9�r�O�6�о
pܺ���0JN����m�1滃�������;����s��G��;	�F��j�E�����<UƱ�.l Wv ;�|#�����B�/R^��P���E$<�䝧e_.b�ڸ�����V��sf�0ʳ�cߗ��U�"�X�9$�Ob(�N���T�1AgR�@�n����w��B��v��\�X�pZQ5F[k�D�-�s��W�MsS&g_&$_���3�}i�g�or,3�f��p�]ג}��|$��2Fɷ��R]B���c��hn��\Êd���c���0BT�^;�f����H[��~
:^�/ƶֳ�q����ٷ�vv��6�[���
��$5M.�k�[7<Ԕ
�!0�[���k�	�C8Ꙣ�4Ia��җ����wy���]������vI�tZ�p��"oi[��3 +ذmO"�A㤺�ׯ��l}d��F�"�|M�ulC9%+�0�Nv2�+��!=�����8�q�R�}P��W�9�m}��&z��ĉoR�C D.�kD|��*������ZRxS3��rs]֟�	�s ���(�=E3W3�T�1|C);)TEv�u���s�D�d��K&z�7L��A�U��y����u����ZJ���B!��:��SZ˦S��6�&֩���]�K����h;�^Xd����d�i]�j�����7Cyf�ON��K����^�J������}�G.�lYQ`1;ai�M�b����H��>85rД&��Q��E��"����a����Ä�
�u�i�^B�^6nR�E��W NXۑ�R��h	�Eɋ���-S���0�[���b 0���j��7���5�n�/��٫ݵf�T���"v���5��b`g��{�k�v!�Z�6��v	N,�As���Xtc�5W	�^��A�m�~%[���O@L���[����#\�������sՆ��S����9{�B�����`?p$�S��=<�;@zD���'�����3��B��[n�k�^�	�d�KAP�$Z��H����k��Ƽ	�N�fF/�h�������%�r�?���.8w�(A���\$S8b�9�Ǟ�x���W,-�ˈ���W��ow\s��4O�YV��MR,bI@oϺeѭB�;�FY�z�@���#֛�nٵQ���Ld� =�8w`R���[~sڹ:�1j���]�A��*-��x����q�?H�{G�s�}=ם���T���ڥ0?X��]�J�'�^I$�̿m�EBQc��帓j���_�Yڐ3�f��������U�X�s+��R_�.xg�����Y���[�>����?xmlJ�Bߝ!:������߷��4���d��#���8W,������C��cc����1iu=�|��m`�ܼ��Jy=���w���#�u	{7Ub�A�B�5�jd|��K_�����*1�s�M��%��d'-�\�5bC�J�����F@?�ӌ��-��@8=��9�(U�`��h��r�VD�D�˟�xMqd�Ĉw����5c���������U D:͓�����w�h�n���O�*hW�P&�>盍>��|�W��RZ<�	���m�\�y۽?^�5A�{��䟾��w+�O4���į-�e�T��_���$a�ys-I!}�Y����Bm��I0�Bag��;Gr�qٵ�C�x��0��ֿ�����v���3H� %L^JF6��9��<�gلKqKT\��`�t���k�������>�ە�Ao��v���𙱁�֏�l&ܹ�X����� gQ�X�?]�39�̴x�+A��s;����[��Q����QQU�W�Ȁ6�5}��?9(�
޳��	)�{�'���[�Tm?�Rf,E^�z�|��;�|1�x��~�?�� /�e}%�
W�T�g�ɱ�O3^��Fb���F(���WB����-,��Ai��S�Sέ~������w�P!z��� �Z`?���� n�D|�A�\�\�Jv�~n�)2�j�3����و�DH�<�\�\V�q�;���~�^����J��M��>g�{1nlx?�>�ߞt��᳉j:i�'o����2rX���XHC�j��R5��> (����1����8��?\
Uj��}o��8��(��eF	e����/���Hs�wa�TS���ˠ<gx�28Ο�>CaB���N�f���~�cl�2��^H�>@ht(Xc������!�c���l2��9���s���;k偆刡J[+����M~*������'$_�T���S�����[~,w�7�h$C �8�G��y��2Τ޲��e�����-�A��Ap��,��2����w^	�F,?u���x��D6;88g������k��3U�-��I���l�N
RӺ�c�.9�nx��E�D�2'zB�}u���y��
�w�OJ�m���\��o�
�mq���V1X!���B�h ��}��t���k�
ҘK� �.��ӷG6�s�+�W��Ŭ�i�u�*/U��H�"h�o��c2�{��|b�#c�4~P:��TX�8S���_��k��S8�W�b-�<�WS�Z�z��k��T��B<�wN�FH�P���hA����'���x6:�?]�]9M�YW\n�l��Pi�4��D�$53��)�!��#�����y;wE�Q]O��O�mx�:PT�	Bn��C
�L�	�,�q"m��������`:0t���*?��RƥO��R�'J�ڤ���Q�*>%f�wcR���XoB(�;����t�^�|��b���k[j٨��T�]�ڂXÄHn~�q4�x�-ۛ�(��҅�&^�8��~�*U�d{�:�`)��r�"�o��#�2
�h��sDKw���Gd �@�\[*�\�5 l�?c���l��{�+����5r��1��Θ����40H��}�m��e��:����{*q���@�=啔���8x27�ො=6>�=a牫ԓ���;?�C�vN��ھ��>��L�}?��IcҚ
��y�-�fFH��Z_c��2�)�~7�>mЙ�� VT� �x�Ն�v""W�/��?�h+���')�m��Ȃ��5l�;��G��#r�H���X=��`w�@�`bևet"9��\�p;rF��d�����{�Pu?�_��&.�8&�$�oEM\�����cS~�6���5#��Y5����k�e갟�� =gޥ����4{��/��͢���*!���*��G/	DJ�S�NE}������оi��V���N�b!�fodW�,&u���*�i�4�����\�k_��kr�܇DJ��>b��9�f�s\���GdFqC�+ߖ�W��R��Ħw:f�>g}ݒ)b���-U��7�k�=�mz\Q�.EIS��Ţl��oN�ws�܅xLH��[Jb����l�9i֦�A�Lc7�P�Z��<������۩X���w���c��%�����ڋ��y	Ŭ;B"-�.��y}��ƹ�fˌ!�p(z_�Qآ*���y�6�U�@ a/�2�q�ζ�li�}����>܅�L��.g���"=:�m�r�D��K=�@kD{�#�O�l	9�'�uWg�z�W���G3�4�D�f{�kﴁ/�U�t#0&?�{�2ENv���޷	�;#�۱�����$(�q��sL,�f����.�?Z�����l�Hݏ]�����O�6��N�2w	.1/М�7�v��9Rt�W$Ĳ�Uǉ�/�K�A�XG:���]H���k �g����N�lK%�o!�Y����)�U(�I�9�c��4��z>an{ ���?^��y`H��91_�o��#�fd�j/�h(�P\�<ˎcM��@��1�d�i[�^�0ʞ����M8�����ޮ�4[��1K�W��m�u��bh��wVV(y.�y�9syp�< ��}h���c�u��m8V>�AT�_7�M7����jl[�;���'����\T/�����RM��?3>�ӆ����*p����й�I�*����W"LT��H���\c�_����V>l0<F�/�"��j 8!�ѩ�y������C2��`��JJ������Ʃs�{�w�G��)I:F�>�f���9Y�D�ӉX�aH��������;μ3��3o���$�����&u4�P<p⎃j���x�tKx(Nf�KT�WH�
�MW㑳�p%>��>� Z���� �ܐE�c.��0PߣqFɎgU�z6�ɗ�g2�˧�	�d^�{W�o8*���km㲆�̆�"Q����?'�-��<k��3�����ݻ��S���pF�+l.�ю%��T@MN7.	�fì���9~�d-a� �y{a���){����8[�S+����C@�M�JP$��΄��܎b9J�D �2VN����ut0��_�����6�d�^�W��ݟ�f���%�NДu��vGZ�W���$c;�G�RZ -���gm�8�cb�g`~���'����"��Kb4WlA&����:
:���x0�h�g��0.�(�BqG��ꑟ����&�I��ȃ��[��>;ꣾ����|�<�qL�Iε�'�#�K�<���)8��\����H���W���e1=�l+�~9�e�:�K��P'f��tL��/l�j�-4hA�wxcR����r�֬����w�����ЪPˆk��Gq�3>�I �	���#"�ٹ����q�J�v���町ou&�n��h����J�\N�,a,�x\T���2�{�6�n؄`n�k���$-mdS�1aó�:�N�%fϲ����2��h�N�x�����AӔ�-,����=6�η�Q������{�ƞ���"�M���)H�����O�rq''l�F��	%ZfL��X��K�T،H��p��?f��L���m�?m��A�wT�铵��X��0wu�C�F�	��5�_�6H�J]��������<��'$���Fqa4]	�C����	V �w!�����*+k o�&�u0��:�)�uW2*of�*KO>K��6x2=J��&���HU{�\�63y+#8�G��h�)-��H��N���(�r��`H�$�|:��~��T��7�����L��W-��`q�K�Ʈ�Fo�&;=1[U�5�?j��.-.�z��A+,.x�o1}��n�