XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��/��f���G��츨����_۲�5��6*����Bu-ً�LC��i6b!X�_g�1S��PP��#�EY�V���<�YS�|��jz��o�˓n�#�b���ݒ�z��-="��>0�|�]�-��H�IKf��v�[�'M���qnas��abֿP�Z�KC׊���[s����a��pvỼQ�6Pj ��r���gefl�[-s���#�6���)��@H:U���B>(��X�^��K-P�*��NB���U<t�/`��/`s*��:����z+r�I�v�ܒC���j���IԷh���K@:3i��{��9��~&E�mw�]�Z�V��wX{-쬚�&D�C��d��՘7NE2�1��w��A��8�vG���Qc<�D�� �(9�/T6������ fs\��n��va+��]��s� '��=�oVEB��Io��aD`װ-�i٣�� ��V��I�ѧx_*�����B���ޙ��#ŊL���LQ�^��B{�[�5�f�/��vi{��GZ�����?��u�?��L%���G+H"���҄%�'��C����)�)���y���8���=D�0���{w5��#Zu {��`�KXǦU8�\�j�YrlR�S�ד�:��ΤA�c�4,�cķ}n�H��7�\�2G#��vd�d˃�R�%m��"�I*�X��eIO�)�g�f<d����V�ߨ�zV��+z1�ԩ.Q��Ȏ��8���ZZ�����d���+9z�)u�aSW�XlxVHYEB    fa00    2230՝1�����f�[��N�2�i�{-�`R���zĎ|W<˭�+����:Ogq����2�DО��5��[k�Q .̆D�u�"<�9���j�����:����%��ȠXu>+�)�D��(~�!��H�[���:���j5G��Q�	�f��|L��	�_eEt]�<eގ�[nֲ�^J/��S��O܍K���K�fyÙs�y�3�?�Qȗ�&X�$����&�#\9�x5m����j	o�a�I����7L:� ����_	�í:��J�f�䵊#�����:��nf.�p�KU�?%a^�NF2��m�������)����k�� d�IZʑ#��!բLANso�[�o�ͧ`>Z=�OB	�z�zm�K���Э��{3JNJ��_���\��䪞E�â6(S&��ްl^<T}�8�Н����'ډR*��	�S��
ĸ��@V�Ly,�2�TZ}Ha�_}�N��;���[�n"�g�*�#C�b1�%�E� e��z#�E�>��+���Se[����PZZ�mxc����n~D��2ȳE������rg�ՐD\�%�Bq�U ���7E�{�^�p� �?��͞ߒ�� �&�TO�Fm�?z2�H`D���]��w��`�x�`��,La�.�����U�H �qFw�_ e1�f���U2����#��"��v�$r�#�4��937�;��t.Fh�d���̧��(�)��+(EѠ����x2?&b�҃�8Y�F��r۔��}T��֢3�o�]c����}�OǛl5@�|t��ޙI�T�0ZRmã�u��%X|UDpw�&i�%6��Ͳ-�f�`j�ۉ}�Ũ����,k�]E��5��K��|P�"���ڝ;zUN)���ȞD�Jn��Pл�5���xGb���q�5f�D�.��e���N�M�N����.V���0���#�y_�clH��;��M9482E���1�3f^����m��s��^Ǎ1�{����o�*Ò���WI���l5�h�*����YJw�9Ÿ(X?ℲTS��k*�MZ<����=�<Z�������1ϣ��zd�`���s3<d?����@yj����a�uHў���̇�G�~��o�>�"�k���׊b�c sh`��@��>�,X�B���(�.���7�ߟ�����׬\����W��wĩ�uڍ|t�X�	^�)�{:�0�s�qZ�H,n�*ȉ��ʦN+�e1"�ův�;??����zZ���9,<�ܵFgh�7�k�V7�s݅Y�ߞ�L�:	N���|�*g���Q�i���@(�>ӄ��࡙�� �	r�#���`�X��
���Vbb<������?v.�mFĬ\/��A�>`��^�	\�<~o�+Q���Zs�o�����H�"�� ����\{$*�4���mN�jl�ތ^�
�1��C?#|�=U�|���������� ��Q��W�K���il~�OƧ��E1��j���`2]1ӧ�Ѽ��!���s�~��X�754��͟&�'��M68��gǄ3���xd"�X��/[CV�^�ʂ�a��VK �J���t��A�����&ʀ�\�����9&��[x�`��1��/o}�ef����U���� <��tHG��Z�0��m����-1�`��}}0/�XqZL�4��w�`]?Rl������Щ������#psYftr��:�d��k�觩�f��-�N�0���c�?� zo�xOP�G�TN���Z��=G*�q��z�t��X�\�����t��l���|)^�_�ip��ơ̇����:�:�Q���P�!���]����w�7(�a�(���0o�\�Œ-$�bdb_$~_{��"��#�į�Ȋ��A����s�6K�q~!?�UDkt���D�U ��Z�&�07Ad�i>�7H�[j����k�8������z|l�^��#p!�Y��o���c[���3���+?����F �L3��OE�l�����أ���Ŋ[��z[�b+�5�r�"�cd��yҾ��I@k��^���_3��	e%%<�򀱳]������"^����&h(�8�`?ɿ�̞�Bt<�,�� ���;�C%����b�K��~#�5[���g�sާ(ou0p5t�7fܻIr�TIwUs��|�ܖ/� 6����i��z��,���]%�C :�5;�"u�`o�m~�t�?Ա�����7	^$���Pl'�e�"�U��9@�Y)�<�3��.&H�����Y�_b�ӈ�@ܢb;R x�*���C�v�rX�!���֠���fpS��w��b���,�T��T��i-�$���gɉ�<P�;#f8ͧ��mx,���҄�o�E:%u��'F���C�vJ�8PB��V��E�I�n|��3]�%e���ݟ�-�Y�C/$ �����}��~��������&
�d*�n�*��Eۼ=��2����4ko6�G�-G!�3�;c
���`��τ8��ǿu� �a���ESf��)�"��j6�-�~�9��1�o�ʹUuU��s�]Z{����r	���#�sh��}ߞ��9���|�k-y*�
gN+W������^1�4P�Qd�m�_���y�nT������c�ť؍ ���I,@��
�<ED�Da�K������^ef�����:\��N�"f̪��X��<C�vቶ�;ɛp�nM{�/�!��;�w�%,`�w����� �:B���#/�����w^Ǉr�M�S���I���u(�f�j-�m`���$�or�Q�����	�wXB��,�h�d���a;	1o�Q�c:��qj5|�U��.\�Bwj66��ɏ��d��Z�R1�PO�-������_a/�(��dA�����6�Z�_2ii닩ڃ��ʶ/���V���g��Gjk�O�E��9<G�.��D���<��/-������Pg�ޫ�qX�ʴ��u�H���Yk�N���[��z}f*-U��sG&�U��`�~�|`P1� ��kN�vUϾ�u�w���o�U�8����)����:�Q)�R�`e�#т������A(>���Ǥc�ݾ-L�>ZG�i���RJTR�aN�KǱ1
}��|��q��\��t����/O�;HU��Z���z�A'���Z�	�1�Ƅ�����`���W���<oB�o,�[M ٸ��x:2�p�Pȇ ����\O�N�Ҿ�����[��3���- �Q�w^� 6�CҶ���G)w2�[;ޟ��]-*��H�����R(���t<6-;p!h�w�)Esc~̞;��{:N��TEki�D�w�X��?��o�}��� J�A��Ǫ&a��:�0��TH����&�p�'��5�Q�F&cG-ہ�ni�;�{:���#�Vt}��=��1D.��_�ɟ��5��)`����F�09�R)�Ϛ�I�`_I����zwԦ ��|���L4��ʛY��0�D^
C�q��":;��c\�h(v9&2j�ˠig'��o>w���°��(R(7�k���v�C&"�(�7��&�V)��p��C�ųKW7���R_d)�c&�=�u���#^j�9��񾈡Pf��z��9(C�t���{1�o F�p�b���Q'���e/.|����2���[/����ι���/����ʺ�$��$����V8��H��x
�C])$ڿC!.h��x�}�v4�)M��ߡ� ����������[D�ǹ��4��p9�RS�|�.fL�}�!�`!���'<�"}��9,M&���E���������V��A�m`hd�:l�������ksA[UrBړZ	E�s��lO8`lt:.����gY��,�6Q[��S=�ˇ�Qz��jK������Tx�PI~P\f�p�|�����]��i�"�/�ő:��fk�P�S3(c�Ud=~��e�ګ8�2��J�����`a�y{�z��W���:�^��MlLoD�<�aJ���J4�PS�c��py�^��>���{E������!?P��?h�����_=�S�ڶ�����	#]]2$�D&���g�ֲ�F'�>�s�3LV��OW�`�k`�P˳�ld�꧍��S޺$�����5x��6�	���N����1	B���h��ц/���[�q<
=$��~{���_�p*-���.΃��\�W����0��� �޲V��ό��Jr6K���z��s�h��,�Z�l��Di�1�E#�[����:�.�TU����]M��"�z�@w
��IV���T�K2�^�0�d�	,��s`ӫ!��_OO�'��N���Ю��N��&�����gw�{�A�}��n+��*Xs�<~��B�C���1�gN�g�e�]�|�U�K��7��}�B��,I�!�@=
��[�De� ��;p6�9fWڻ�t��4��;�Ņ@���ϯ"�������M���i=��+��Əǔ���av�J86::�h��I�s�~%AC�/,h(p��X#?�=P��b1��}�׀��C���Y��?'ǈ�
z��EN��c�a&�̎��<�ah�:�0����0_+�|�)��-]ɉ��g��%0��7g�2o\9��AA��c0MG�%�l-����3�}�����ub����扦�ˆ����ʠ��%e�Fc�K����̠����B�Q�J�G���6J��@"Ff�:�Z-��|�g����;t�~p>��7ELY��o�������7��c�����~�����e�.nL�߁�����"e;�_�����	TRKKetS��g�d�AZ8�����n7��9�C���`҇��+�N�F�'v������o>����!��]2�oA��^jKC�\����:��m	։S�������%��lE�g��`�<��៴#�T�7���Ǖ�ws�tH�� ��;t�Ы\|�<!w��	��ݫ��v��t����U�?F�|ƨ����W�1N�����t��?��t}����� k�T�)��������f�:����M�U�|s4���_���j�<z�٠V�/J㜬����z2���R�1��8m�)u���U⦏��݃)N��@��d�C���N�LGh%n����$�s~u�I�-�?����@���G%u+����.�@�#�9�~�=�tW�]�l���$| �Z��zFE
c$x�DF,�đ���`�����v���P�7⤎��z.��,#,?c�j۠H�;hk/m����ҲD�������9 ����e����"V��J�"SIJ�>��+SK�8n#̐�?�8��{z���ʓ����*$��6�x�oQ�[�ܠ��B�@<�u����-��z��b�Bs���"�˳�B]��=!H���J�e���7>��T\I���ӿ�C=�x�S�<��K�	oW�&�=)����I�%D���z-��5��aQ�л���qGb��`Q���G_�����Z��� ���< �{���E, ��b����"FEC������`�z4�I}���%�7��_?������u=I���L�$	/��*ٌ�W݈�>�-��L'6֝P�MĹ�1y�Y��Ls�I�u_�<!�#�|W(N��e�:���x�fx���
��BҒ�d�\UIWߎ�P�kr+$nֻ�ӈ�{ɓ.~˺���;?���X���֫���Ǳ)��?I'W�kq��6����p@P}O�Zb�9m%o�ċ����cYm�*x�52��|��u�Ddp��$oQ^z"{��P��=W�2�1�l-�<5ńO*
+ne�j�9�	�&Q�O��HoJLRD�\�&�y-N9⦉9��$}���Cuj(��z�m��biA����P��Κ�>���{����ߐ�4d��2e�a���a��*��c[o%)�Qס��k.��yaJ���	�bsf�w%tZ���L�Z/�2ȥXe��j���H�iF��U��l(餖(z��$��j��ӥ�a������Q�f�?�}��~�}:�GR�qr�u@n��mY��\@��91�N�-�U����>���{����vR������?���5r�!	�>Ͽb�sb��G^��su�tR����ی	���\��˿k�����,�Fl�����1���p�<�<k�۩6��*L����kk�A�ٹ%��J��u��U[o���=_�!�d����}x!���o%�U)X�k�����S7�U�șS��) т���:�{�y��d�.^��-�O8�cF'��ݒ��C����k�Qy|C��.����z�v��?!
�f�@���h��su��U�@W��@A5�0��е�`<�B�aZ���;$�rA�?�����M5We���G�
��(�4���HT�i/�r�7���.k8�؝����uЅ��K��M�Õr�^@X�g0��I�y��M�""k��wj���o6�:	�s#�~�}��.}'!�����L;R�h�~E �X��=iy��;U��'���?ڜ�*O����.}n�Z@A�m���0��ʜo.��"�d�t�qm]u�{d��0�w�7-���wh����)Y';�t:�p&��\�2�{&����a�g����b{+A�fB��Y�M�Zr��g�9P{�!�d����<*����2���|���u�9L��U��YKm&>34;����&�
o�MZq�Wc~MՕWp����0s��2K|�'�Dd�:X�� "��M�/j���D҅{�~܇�}�����׌��G-���*�$\���ވ9��d��]�'Q�Ĝ�yh�/�y>$�+��O�
�j��j���V<�B���k^K�A� h�;rc9���;�<K��+�Q���A�A�^�@)i�i ���N���Z�֤�!� �r�?R6�S3�����(���Y&K@p�Xq�vݶ%������$�X�	p1&�!p�'-:f�0�2}��ñA���f�*����v
��̪n0��,z��a&sg�r ��؆6�h_���7@���%|��v�0����[��
�4u~܈f3bn��=�7ؖj����N6�Uܢ"b��3�����Q���ަ���~��m�����_hF�O�����0/N���y��pEˌ�`�K!�'�ݶ�3���8&aqpx|���әGv�U�OBnw�;�a��4�6zX�����M��h��	<���
 �pvÜ	��7��2
�,)x��'Zd��|��d�Z���,�Y���������!`NՠS>�x�U�^"���CѺa�b���O]J��9�ȍ����1��>�vdǉ,����^�"N�W�����A%sN��2��-P���_B��P�����"w2<����#��s�?1�*��R���򃕥��϶|�jr�[�.��z�zo He2�י��}Ձ�2ωq��nG�sHM,�1@�X���y�a���si]>	�"��a�����s��^�%g�>��wu��T���ַz9�Џ�V��%v��#$9B�*�-�1����- ��n�U�̷Q�7,�.5�&�sF{��Ͳ�t�Q�����p��G�N �'��(E��D�ޡ�����`�RI�'|2➄��3��8��}�3�mk=$ħ�fZK8K��u�s�h�2Ȁh��*���A �]�z1�m[�)�����suk���glD�k���{�Op���ϧ��C�O�c��l}kmkM��������f����YvV��h��: :Ʒ���D�|Px5�@{�����Z�A���"_��;�9yt� Й�I�H�g���{��c^7��jF�1
U���ߧ-yi��٨�	�]+"�����
#��l=5�ĥrA�
��5���W�1%nCCa�GR�<��"��X���v��Prc�ٓfJW�U�6����:Rx�P�k�꾧«-䝰I����!�'�ܤ�Ϗ�Lj.c*�I��KɆ�Z���b.J���/�]�� ]�ClA�ǉwa2ܕs55:�WҪ��N{H�^����)ʑ�z��-��w6.T^��������ա~�C�:T�<\<Gk��p��7�n6i���k7��숃 �֒�����,��!��P��z���Q�*�Lݚ䏖�6%���b���j:x@�~	��LAi�+z����\����p�GB�����ꦖq��$�9��觚�1uM�����!E�}k)���7�{ֱ�Q0J]��G�Ĉ8),�¦�,�K�X�W�N|�̴�VǯZ©���ŏ���=��@�v! �Y=O����{I�#;>A9e�0���J��p�*��כ^��=���sy�Z�M�S��#����aⴻ�PW��ܐa;q�����d�Ä���%E�gRg9!�G3\�Q�%1F�S���nR'CТ���v����!)��|��3sf���g�����2Žif@�����^��?����*��c���]>q��=�Q����Z�a�^�e9��}�N�H��ygZ=����Hw6�$�!׶�|�(���ddL�,˦��(�X��Qii%�R��᥵1nw�)�*Z�%0���.�S�!��>$i�_�E���b�/�K�j�Pc@�˯5��(�4�-���P x���;Z�����!9�4B�5.`6�.YR�r�F� _�Dw0���`bƸ��\:u�l����w�߻�@c�hXlxVHYEB    6682     5d0$�ۜI A1���Z^�變P
ܙ�R���|)-m��{w�Gt��A6���+=�t�Ӣ��$(X9i����/je����Sq�MZ�:���߸�&?Mݓ�?�zJ����Jo��~�G���1a�����=6�`����l\޾MW�k���a�p�_�S)#��,��l���r��8��G�d���7��l�70C��'#^Q{�2�Q�a��\��E];� �PZA�P?��-��`�*"���7��AI�e���ک�*��MU���<�P��<~������L�G�=,D ̬<j\F���H$���O��љ)��9c����:~ų:�B�Y�
\��5��BU���ԏ��^O��˟
d��@O6����m@>�ڭ]�X�g7�n��ԒHf<�RW����I�h�=�~����1 SM!�5���1�+�Y`���Ҕ�V�z�
W��Ӈ��鮻2��Ob��LŅ��Ty]�#�G�|�5��E�Y~����Jx��Z�&e��0��Ȓ�a�̧�L�r��}����q;�]���3�Ep��(�S�j�uiU�ܹ9�����
�~�5�����3�s�V
���:6#S�i\	���$�|/�/V�`��ݷ�)O��8P,�&��[���t���͵�k۷��׉]�����uGI(;�	֮�x�m���V�R+�Bt�#��8�|�U�x����D�Ϫq�B�o�9�Ƽ%�;-����K\�K���>!6گ*ڽ���Im�R����<:�A'�D�σ���S��۷�`�F�#AP�-'��g+�(�7��㣁{��������T�X(`�}RՓ_���(�0t��A�1Pl��|�P �E��2�AC�*���LV`�v�X̎�OG
�����ކ>�Ƴ���Ī��;��j�S*RT�i[)�A{ؘ��6WYo�/Gs�%�b�X�%�;�x`DrB}����It��z8W�_�
S\�ʑ
v��(I�uQA��bYƁ��&so������c7ſ����%y�����,.	ݯI�ntA���Ĕ�Jmb�aV���D�I�+ZMſ�H@i�=��C�a�냛8���i��U��o�.Os�Z��%�I���X,��Y�]�@D�o�6�/�yG�j"��SS(1�V1�eV)��TQ�Q]J7��n��i���tbq���_c�;�)mF�NZ���1j��O��W�۹���Ng$&�1��&u�^j��o�u�16aԢ@C�����n��7w:�E��#��2��9��EQ!�� Z3νg�Y��9���=�	 GZ��A��[ũ_�;D	����O������F��hX����t>�f�
4���$��}?\����ĕG5VUԺ�2�h���k��7�
7c�r-�SǃZ�~Iɀa��d�
�8x���;&Ҭ�U�_���s6n���˰I}�"�"��tJ���Z��{zt����K7;;�5�ڝ��������