XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���]ɤ�<v�"��\6�P���u�I_na�
�����#��%��G��ID⫤�yΏ°u��i�Q���=��Ȑ?��Q��on��;����~C���7��%���BqQ�JϺ8�o$AM����i��,�O���j����^+�YM�����l���d��؝����J&��H���+~lGK^�W���	��)1ߔ�B:�⛏����i(�R{���f��ȧ��oL�3�Ep<LW �B젢�ͅP;��Sp��*v�ސw`.�� hI�^��8��eG;����a>�]e��;Zk�"O��K��Jtu�	O��{P`~+��i[��Y���2]�P�E�r��ڣ�ed��ź%��Q�9b�U/���%�p�s* ��)�����^������!ϡ�u:t9J��:LJf,��(���g.��Uic֣��� }�^�����뱮��xV��k�w���EsA�TTo�bp��B�N�D-�S��w��3�F�!�{NY HL<�]Lw��E�����W�I�[��c�����8,��1�� �pVN��w�	��MŊժ7��eCe�@u��1~���>�����5���̃�;���-.�*_;�f��`+�ʢGZ�!
�O	`J�r�O��Z'쫘��3��l#��SJ����):�CR~Խ��!/�-YLc/x���bmg5��Zy?� x��h��j��Ħ���/δ�����hPQ�hY�Io�*���x�>O�Re30��<��5�i�p~�����U>XlxVHYEB    2e20     b40�)�<����k��Yi\�;����k���M�V��� �!2"����G�1~£|@���^�4�gϸX5����T�h8^ʜ�.�ڟH'��{О����~f͙[��R��o��d�u�����-x��WH3���e:��B�;˻w Aޭ�U���fe%\�����
�'��^��^5h���5��\����<���=��!�<D�E�z%�]O�n�b��?�'�13o&ݹx�9E�Z�u����B���s(�w?����a�j��ۯ�X�[c�kȭ�>=Rb��)ۡ랍��S��W�{���R�����h�� =0� e<�x�����|�`9a �:�]��xb��>Ӆ|�惧���l�G/��.Bo8�7���L⧥�?��})�+��bЧP������<����@t%VY�j^��?��*]��E`�(@�g*mC�X����{�<G���G�ˬ�����\]7n���(��X���c)Ϊ��� �:T,�Q��n�$�Q�VK˝�"MW���Ư��|�	��#��m����(����Z�L7�$�i������7곙XqK��,#|t���ND�y��+�'�XL��|BS��]��E��e��*ҟ5]��_�8�T�L�'|�n���Bo`���dex��/
Ę�Vs�n��!x�eK�`i0��n�����ٰ���Ӭp�f�.��`��� C2|*��2�S�
�
���/ٺ�D�7�uqq.lb�Q�n���;9� �駅&/����t�f`����cN�{��77�w�V�`t����,xiGQ�NP��>-�`g�2K��=���ܢ��i�m�W ������0������%�I}��KhW
��A\#�0�a���U�R�a`i囿��������c ���iJ��i�K��s��y=B�R��"dL��0����G�����3�.�ax p\��.�IϏ����%N��Ƶ3�	H���x��$�l"����B��]�i�)
�y���Y�>��N.�H'�ʎ$�QԳ��3�O���,�e�r|h�m�H��^E>JJ���WUKr�F�=�W���t�'>�����  �E�zM�t��cs� �C㪭�?���Il�C��^����.�T�m��[�,� ө���(?�U���U�}vX����߷��	����7T<�16b��6��sBʖis�*�	�V�.7j�O����L�6�s�z��s�dQ�~�,4�t�����U��g�>s�͖���7{T��d�ͩOF�p���@G�g��3���ܪ����qЩ�No	'��mv/b2T���`H��rOy���F^?���
��_Z���(m�ynb+'6�F����Óvva
�G܁/b��@E�'!�-c�w�Uw؏�әx�6o��󲃹N�q��0d<��U�,�����ѝĜ�ڨ�"9�L�W	bA��/���`���8t��������������/��Aҽm�)R��A1{j���t__�21���5S�Ϲk���d�m�wp�76W#E�;�R���Y��`C���
�PD�������ƎN �h�&� ��V���dG�����0:��ʁJF�,7�H]UbbHM�]
w��ZqH��U�J�	-~/�&5QԴ��{BY��ge�d�9nMT�Cʊ��v������X�l[ !�Ǯ�G��E�$�s�S�?:�D��C�!����d����Dk'[��qwEn2vɥ��h"���/8/��L�0Z:�2������%��������{w��++rG�L���@"���P�R����LOT5/�N�I��Ż�?��ym'�)\��'Uj$�Lw��;
@���*_��'~�%�->���qp;@�&@D�1k$�T��c��SR�Ml�n�ԭ]91	�ˏ�G��|��d|&�����1z&	�s�V�^y�	�����L }v%Cw������r(�!��-�K(Zj��Kc�����3�:�y���T�A Bt��km���g2��6С�f����d��!�n|�ʘ�QV�_�9�QR�6��Eٴ�E�'��F���,��х����k��(E�X���e�Rx%��y<��E��Z�W�ۄ��@�"-h-�� �]A<���P��yv�����-�-���*[�Ei��"�����EW��"%���Lka�:i6�03�M.�3tJP�p^�:���2d�\�/3`jeq�S�_��Q����<V�wD�B[`V����)� �z<�v�*��b,���-3�3@�G�i�� X[��5z�s�p��be7g�Q�v��a�:gp.��bXl�wx�ګV����3H~��F2:܄ů�kQ��aD�X��e������Y�#�ad��Jq�(z��(�t?���fr�����`,qijV��I��g'Z���,%�Y^2�d)���.� ם��I��"�}72%�F\C�"%��W>c�YU5g^6:wM�`��)�{d��T��rRz�� �l��!(n�]��eR�x{�y�����6̗����eOΏ:��+�5�G!��5Yr�f)��ԃy6t�����B��	³|~�|&/�<�|ɤ�*Q�,��07@f:�ZyGt��{�f�Mʂ��95h�lGϔ���y��"�q�@���z;�<U����GW�k!���c\k.�#�g���W�#�gd�*��Y�o�k�j%$�?z��q�Z�%����E�Ё5)&bISn�L��>�D�n�a�s	�Y�	~;���m!�MX�ų��`��8�OD38&���
i}��w�X����?+��Fw�t7'���ZQb�C���g��6X���~ly=kr$6I����r �_'�2��N�ԟC\�Z�