XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��5/ɈF5e5��r���;�U.����E>���A��rix���"�D�p,R㲊�U+ƈ
O�[�Wmo�[��i��bb �)AM�C�BE�yꩨ^�f�V5~�=�K�F�~�Q��F���G�P�J��Y-İF1hz�ɿ\�h����������qa\}�
!���$�U��$�RA���,Vw+����
�6�#KR����ۑ�/�H��L���4���KT�XD�KZiI9��ٍ���`�\�=ģ�������Ӻ$ͫ��9�^� ��J�G�.�,�M��l]��d!�����7k��i��ka�ڈ�)�]�?�+c�g�C� ��9Q�R���+�T����V�	����Whb�{�,���	峃������}��$����� �reϛ?���%.���[nUʢN����ܓ�
�F��J!�'êd�LYס,'�ږ_�,P}y��?�@�Z9��W�O�t���3 ȸ(���:h�YHTc�0"6�봿�N}���d�|�n��Z�0%�>~5/��x���p��y]M�����z��V�G��R�[���묈u�v��4H<��#�G�cl��ۜ�r&8�� ������\�-~{?fҠ���Ucq���;]2^����� ����L3�U���a��_�x�}�la�-+�JV��S'�E���+:Oi��D��RΛBY�{Bh��/��Xm�ݪ�Pk^��7�W�h����	�u�1G5k�-��Y�Tڪ����D0��O:�*����h&XlxVHYEB    fa00    2480�mz�F'H#O�l���� H�n�=����2pI'�����]�詵7%��� [N$3y崙إp��>Si���3�kkG ����e֭걤9���ϸ��+}W[�4QtE�	sy)��/�D^��m�
�/��.�~aq���,p��7(W~�B��K���2$��(���� ���=wI� �V�N�D�ԯ����}CQCc�e�lb5UE��[�/�k3�yM�pW� ����v-����x�1������لeY�#�Rx~��r�`�w�
�Xw"�ǹELBBȜ�jՇ���2��͕�2	��-�?Ռ��d��Ch�U�E&��@�q�s�p,wPbX홸�:�ʅ:<��$Dal[�c��mƲ�Ʀ)&'8b�1���"``�nk��$"fj1��o�������*��E�"Ӑ���g7,�gr�K�aC3�o�+��]ցV7U�j�Q5��~�3���A��S���ߡ�O�������)(L�DV�����6籣/���bC��-{� �iK�	M��\���E2�Ju� �!B����!�IZ� ��X/��Y 2H�N�U,C�#�����O�j6���r���Ys�]�� �lE������sZ�׉G	nv�������̋�rVL-��:�;{�]2��\-�pO�R�+"~7-�2DSݲ�T�X `�M>������!����d�[x�/�c��G	�4����gB�_�h>TB+(�&6g��j����w����q�"�US�rQ��J!�-ۚ��ӠT�� �J��++��%D��T:k��uF���O�e�q�C�b�1���������/-�ߤ����Md�T��>�i jn�-�/��Cվ>�X�}��}@���a%Ӓ�Ә���^�'�=�6�l�37j!��d�f�S�j��G�k;��O@��M$
_�h_�9-�}��X0�I���0r1�!�Dg���T�gb��� Ȍb1���
�Z�ku�Xt_��q�:�E�t=Z�O�y�(/i����M&��3���X�-�mB�\��ܗ#���*9|S&�8�&2�0�($�jN�^�R�L�&@&8��K^���O&X�/%�2.4m�e�H�x�m�{g���1Gg�]7٧v�kL[�R���^_2��]% �h���G�\�����dt�dƣP��v�����8�K���3�zU׺�@�D�oKmLun�f劊Z���Z=�o�����Lb�K^������C�;y;w�U�BN�����'�P�c�p	���ᴵv�x�| �$��-;
�>�A�3G�����b˶Y0��tcF�A�ƯX�,i�׉`����*��Okc�EN�k�� '^@���<5����,��)/�S��;IPW�ʥ>'���F������C��~9����Z����v�fwapX1Ԉ���n.>�킠	Vl��3H�Ķ���=F-Y(�9ЧꍝNΜ�`��]�0r���PF�Y��r��f��N�O߻��rtC'�5�Tn���~OyR͟���%��^��ۗ��R}?����u��{�2<i٦�M���":˜�3�~���(,�p�b�+�^{:i���#��K>#�U`Q����sV�X���
 `�=�v�Q���F�RZ{qT��g��gN��Df2`�,
�Ǌ3li�^����`w��Q��W3��?�)Z�ǂ�Y�̓���0��S&��@q�P`ή�s^E$9]���QW���5R��!���S���B;��r��Ndz����\���w��*�^s��m��x�um��Jl16�6~��  S�w�/�;��ޠ��TP
�!v���'[�`������DPK�y�ɼ���@*�G*�}��@��d�<A�y`���^]�K�������q�!F~qM�<�'�1���.p.t��~���~�uLh�Ca�j�˾�F���*%VI^+�j�B`6ۏt��²��<I�����l`��	/��`vnk��E0�s�A۪!Ъ���_�XD��t4��T�xБ@�;h\�S٧�&�d7~��|Y�F5�݌�yJ��b�)���o^�,��c�L��g��݋x�?��ԣ��)����<R8_�?n�/?�{�b˗�sؠ4��4]V�����oH��m���taau\��_�ݗm����P�:��{*��GO�v��y�6�x�B��su5)i5D��	v��p��Y�d�W �k�X+��?���T����I�)D�r�>��!�S�A�Iƶ(�ҧz8��6bNS���TP��r���B��.޸}�=f�����W�h�����"�&��(6l���DoĖFl�6���04�2���0�'��t
���Qi*,L0��#xSj�1�uZ8��n��_=PY(d|��7�Aj��F�*��[�F=�VȄ�x���w���q�(v�b��C��A�)���36�8�Ϛ���T�Ɔ�� (Ϩ �O�)�(6�ͳF3?l��Uc��"�{ډ�p�����s�M>�ڍ� �|���ū�w��W��n\��B�z�OAG�s�lÚL��5m� n�y�i�瓍���+h��(���O���~4E�84�[R��u�zܟ��k
��p��(t�5H�7,[���R
�!.��3u���J0���|�Ь��T.L�1��i�e>oR�X���Y�����E	���R�������-��=�:c^Ӥ���;"���?�o/:e���׹�#�M!��kn��P3��'_�]��w����ѵ�a3��8�@|'�4G�F鈏������Ɗ���}��m�_)�0���*0����ː�q5+<��V�M��4u>e�v�q���6�T�T{VQҒJ�	VͳxAc�㕒	����J���yE#��0�*ߠ���w}��X��/�u_7'},?'����E�;i$M���p��k*�:��yt�$'h>X�O����Hm����D�
����q��#y�@bARAS!��5pTNƽ��!�QDFβ��%��$�[����1m���g~��Y��:a'��Mqr��dRڦ'X����_�����䶟�Э����A�e
^++�k�ᤴ���:��&t�W���k��tQ�Q
8,�G�,꺛�����ܖ������y�g�_�E�\�H��c�����ּaۜ"�]��2��}������Q�11>��L��3=
���b8�^�j�Y��Hb� �¸Ux��� C�[�w�H3̿�"Q�Hy�����4�2��ٻ��^�̹�?T�(1������)�wS)��
�"��w�tˀ	D���0o����5�˛�S�y
X�N���۸ �Vd;�����8˸���AD���-�op�.���B�u���%�}4w��O-1�kL ��,*�p��ǚ�̐��ܫ#�>�s�0O�V�-E�J���cM�>;��/�&�*��$���� �HaD~�]|���}�u�<���O���cʣ/C�k:�7f?:jJZ�����$ܞ�OŊُ�S�-y+��.U-fk)+��3a�Y����UizV��z�k	�*�3�N��"h��9#ی"a�ֵ��5bR�z���R�(�g�Nf��^��ܻ���g�o� ��B}��2KP�d
x�3�{���I�#����h��\�&�{�{Vp]v�RehT%��@� G_�5y�"�r��Bx����9Z;��"#.��=@�=�<����gmbeN����7b��ĸ��ρ����T����$��>�W�ՖVC�J�.@�2�.y��P�H�~��\�g�;���{���5�a�k#V�h����/�)9d�]W�7y?=�2"���@�=���JGAM�����{C;�n뷭�?���������4]��{�ѿ?�&	���`Xݱ�uy����B�v���g��� �\���y� m�t�ԃ�*��)���Ro�6XR�*��ԛ+R\��2}H	ż<x\��t�.k��[�y�C*�z�~^
�&�� `1��ⷘ�|����X�	j�� ��՝1�_<�~4�ﵛȡE_e}�Eh<#UF,^|͆�j-�$R=[�8�~0Sގ��lV5�8���6��u�|撱|�Y�2]��N�@�㙅:����f�'�h��G�M�u)p`s=��CTIHR�M	R1v�M=��.m<���� �ډ��a��0u���x;l���vh�<4�hѨ3Fv��FY���hZ0\�Џ�۳�;":Ikr�q�܋S$��t���)T;̝���)������D�޹��	�-�z׵�Djs�ӛa�.�ڠ�L���@%#�
�]җ\	!y���&E7��0*�ل�.=U8����f�[5^H�fp
�X�VwN�@����-�%E�S��G�)=i���RL�KS.�@$;�"=��N���(��!)ۄ[䆬��m�md"�����*Z>��Q�,��/�|4c��҉�b�'[ ���C�X存�+pD��i����>>��V�	��d[E��עC�b�Bf���}�������)
uz" ����vqE�����h����qn�i��/��Pp��և�7���Ң?��r��'jSu�h�x���LA�*�����@U�51X7ۙ��YU!�i4ZD��?Ls��<�Hs=���U#�Cl��P��Q���}B^�� �tX��Voje��������=\29\��Ò? ��4���H�h��&74&D��z�s����vƉ�4�f��2�Imt*MT�K~q��[��^���	rM�ƶ��X�WˡC
.�UY�m����faU�D��A�g�-�-P����.J1y$�
��^8�+]��9r�vu���z_x챩0����} e�G�m�!px�zG�	1�A�<�6_��>7�;���'V�K48���/p�7̌�-��y(j�N�p�!�+���~ί�=I�b$q&�������u��'��+�ˎ
���2��7a&O��Y`�I1I}e�~]��_�uW��&o�$z����ʙ���Bͦj��{�0�'ޞ�ǃ������fw\-�D3��@[	���x��8Ӈ�Or���ʁ��{�(��"]�� ����ٳ?��$���XN�`�wyW�(d���-�Y4��JΦ�u��?XߛHu������h48���Y�?�]���t@�wPe�� {;�/��0���c�{�+n�ظ�;Lf�<�!�J�����|5 ǦK���ݭf�>�{��t�S\T`N��z֮I��Y:w�����
t5̔�ƶ!%�/���piF9h�K(�g�[T �,K�hl˷S�)��3��Q�I�x�u�~V�s��T�p*yT:`��X�L���!�8�� r�Y!��d�2=�/w����#}��+���T�6h��t�r��F֐3�Dc�]߬�"[�aC� 6���u�}�L(R��a8��㺾��uC�W(�xs����f��{�������ai�H"5�[�l[A��~��sP��e�_�6;��F��|V6tv(o$9�iΓ�=�ֳ{J�zb�Xb	F9ʣ���}�M���(@*�*���/�!�$����iH�w�9�Ƥ�ބI���$?���h�H��G�N�������+(��EƠ��ņo �_2�3���x�QѴ���'UU�_����|i�.�۷�n��#�&�ǀ���e����s���#Z͉]���E4]f�]��wھ�+e��^w���UM7}�q��)<.���-��>=��\lD/�"�8�;��̚ꠃ{���]*���A;Sv-c�wn����{��RL�x�j1�	Ԝ�F�̶f�NuU/�a>T�ȸq�ad���:,�K��;B3�;�=d��<n:�plա��s8� x.d�K�x/��E �����m���%P�R�`�u�p����`��.�;���o�b�`,Ǒ�w�����%ڿ4�	���0I�l�7��Q�;�@����K}S�ed2DƆ�ԁ�'H�>h�[�+������Xa,�T�*՜�4 -��Fw	��0�ah.��;<�I��j�%�L�69�0QO�3�߰��@p�vN������]ƪ�	1�D��V7l��9j��G_��S��%��r��'~��^�	o���0��o���/_�w#�ۢ����Z�X����0�gEH���R��S�g��,�@�(�� �Vlk�<� ķB�Ε����:�a�8�3S�^��X~�N��#��[���3��V���g�_ Kń6rae��� �7�`��n?�mW�soPԞ�hr��n<�3�@�j��-��e@���o'�O&�V�Ңdt���/;.��S�8��v�]��J}",��>DW�dWr�G�)������)��<����9�'v��yc̵�q��Hc�>�J$�l�T��^���>��g���+L�Uq��3����8��*�M���L��Ӆi�87F"�tUM�r�
�c��2�x���Ѥϸ`��k=�$%�B����c���nН�w��y"r�?N@72�)��̪0��}@���
9����]DA�!���=q� +M a�K|�ֹ8wvzHuq�_ւE�;�׿��Aݕ�w��G����]������5�k�F����rG�Dk�oU�?�o�g���),�n[�y1��G~�]�S��\6Wݮ��5���dL�3��<_����>Yf��8��q>�bog\f�֩O��Z}������]�M� ����ԃPˣ �V;p��R!�
=����_���.M�Z��`�K^?���pH�1X�w�Y�å��]����O,H����﯑���Q�>�	�IL���^�s􆭽�:�C��pd�	'A�ê���8p�Ա:�)���?�볣���_�a>q�s��0�%~���jKt�;~�S��2��/�~?\:�4{
g��|�{�����4t����@9��vB�/��d��pn��� .��/s��D4�X�@�ۺu�0S�˷�m�n�F^���y5��-�L��J��lUj���	�i�a�E;\���r�9:ޭe�:��)�E���ѽ���E��D�Z0����o0	=X񺿣=ÞQzxNܨF=U	�CHg'��MI*	���<)��r�;=&�u���4����^�E��5��dGX]N��'�T��j~Ft&4���ˉh��n^C��Ê�H�V�5�(���]�3*P�WӠqxC%fޕ&8��A�a�z
��O�Ez���,�O��0��!N���� ��LX%�+��F,�珗��=d/�Ӈ�Ǆy׻+gXY/���c������+��ʦ�4���rP�#>��s#Yk��k�w��d�;F#Xn�dwƃl�%J/h�ʂZ��6Ua{�	�����pO{�?��\|ST�C&�Kg�\?�)0s�*n���&�	������~���� (�%��y�j���J���=���ߣN�Z9�qT}tS:0yAgi���'ȞT��E^'%��I�WT�.ۀ?��s�r���������'�G��^���E%�_���[�h���a�tzru�Ej͘5�@$=���.f��ԁ�#"����nN�Zk��r�m���z�w��$�J�xxE�V^_I�>��{t{W}@?�x��+�ç���#����v������j�O�����E�\�V�Zθ0��}��_|t�5;��f'ٰL�g�M5t8�N
�|A_y��YB��Fq�t�%_f~h1_Ǖ��"�+Bb�����/I�W�~�;8ۘ�"~Ud&�݉���H��h��Iɸ�1�� �&=s��[=�&�a� �k+���]\���'{��{P:��;�+,N�m�e��h���7�����ڹWv�"p�Lc�kj\���j�&���� ��ݹX�Xf��W�W�����K��b凔F0�ͻI�h�)=�>Đw���N��{V)�,�U0���Y��qs��N%�q۾��O�������@��=�?zM�x���Q�s��,�~��嫰�\p��y�kB�E��{vh�ˠ���# �v�u���m*M�94*�f
�R)�Z��1��q�:HXs~di�� ��h� ��D��ҵ�:��5䷩O)(�+�:i�����3��ˢ�KV;@G��K�ݼU��׻���!�\�2"��yr�^"FQunGmwFy6�����Ab>-ݫ��V�Tڐ�h*��eWT�.���w"'�-�(�"�I��#x��r1�P=���J������� ��z}lh��2\AW�F����d<��ic�z$����?(��د�%s�����`��-k����9����i!L�#��E7�H\�CD�'K���-~�+;���2-Ұ@�}�R�A������!W��ѧ�Q��=1@A�؞�����e>uf��8�h�J�f|!�N�YV���ED?��L���;ݸ}���\�\�ڄ�H\���
�<��_��.~�i�o&U�`�w��.0���3|�*�J�I��z��������z�5|�6�w��V#8�z�����M�t��b�����m4�,;���ԳC/F�O���#���^'U4����O�d&]cK7��M,<P�;��m� 66�����+NR0l���h�΢[��jSaʌ��D_�������О�7'�����/<�yd���E�����)�D��=����6�%C�6,ߦ�F��7V_��$��9�M�%T�ږ?`F���yx��?���y��4_Bx�P[Gɔ�!}n��u�#��`�gܳt�0Q�׸���`�6
�?|d�ה0	�P��b���u���@���eK^�����=���	���WB�D����֎F��q�]C||6Z�� �\�.���E:��A�GΰH�8��#-N'8��b���ޮJw\m��c~���������o?D��z���YٗMX)���L!���öfz��r�p�eϺ���1�E'@���)N��ʪ�΋�ä,���̓8�!�u�,���{R���0Qc���5�+U� ����
5����g��ۢ���������Y
�q��-�_���(p�� ����@�v�[$͐q��hY!��ˋ�ax�6��~��9�2�r��N�:��^"c��Iÿ?8꺷��H
�����'n��5��Z��Ӡ7◟9lQ0��lD���f�K��c�ZZe��[j��	����Օ' ��t���D���r>:�oY_��A���Ӄ��q�~�ݵ��Wad���L |����%m���
���1�P���?�?�}XlxVHYEB    964e    1150��/B�&p��P���Ly��_k7�p�8r�]��TP\h�;r�l�d����y���w9bDs[�6�@c�;��~@%)Y�򷙣�K��2�j�{ڒ%B�x�A��O���������tr:��+��.Qn�H�a����h�ߨ�M`�]�(��N_�|lx��%�u4���g�2�2c�2nMNL>�QB�o�Y�J/��q��u��;Z,��`c�L�9�c�G�:8���R��LU-N�oa�v������i�.� �<��#_-�ͅ!�����yK��[����r�Bv�ͷ���x$<Gҏ�����(B���_{�1^d��mXƐ{�����G��%��]�pMx�+(��u&-�~Du��cx[/�W�LjTo5��A�ά0۫��Q9�K9FU����>��%��#��O�x�6����K�M=@iU�]����� (nw�
qO}������Ux�w��,�^-�j����O�`&�S��ڡ�)�BUF]2�K�嗏յx��{Q��d����� �z�i��e*����>��&�=�ݗ��W�3��["j�4:����W,��YlU�:��ӌ��K)�j�o<���}�`��:��$���6�ÿ��gZ]�)�7�4R�q{w^��s}��`�+��T�D���I䠥�9{���ӂL��}�d�"���&]�XM3�6i%kͩа�cp�_����b�'�#��kC�$�
8:�ۦ��C{uL�뻲�l��3����֟�U�9���d����u�]@i�#�����v�x�'N�o��P��ZX1.�Ç���c&!�&)[�t�YD%��ׂ���s�8��ǳ������Y��z�닋Ƹ<��s� q�ب��g�#�0�J��ý�Bjtn�W ��i��m}� ����y��k#ӻ�NM��@�~?8�S��PL=azBs�v(Mx��\��Mu�U�#�FMak#�Z�-�A�Hu��I�@�A-���V�;�Qxz�r��e�ӖK� l�W���}��N�ܛX��-v��V�a>X�dxķ|�h��I���n! �R�'�z{]T�y��Y�/��?�^��mB��4��!�I.?[*�ÁibVJ��R����{�h⹅�X���ځ8���R��ѿ����)�s^A_�Xg���ůQ�d�3�� ��Z�,�e�Y�D}2^[����sT�R�X9uΤ�Z�?�)���"1�_s�nd�����;M/��5��햁j��q�$���y�Y��0��5VIr3q������L���K�)�+�1e������ ��a�W�����XN��ci���:mz^�����{�1���#�S��#���$�b}GҴ)u�;���޼��^
��5+�����3��2u�}�j�Tm� ��v,,բ��fs����]8�Ü��%�K� �r�L<���nP�h{��@D������AMlh�c�Li�^GK7l�䞼+�~��iЅ:f��4P�;eJX|+`&�e�`Иk��xm!QL�Ւ �-ظ®;Č�V���<��u���^�5�aʭ�U܈��+�-� ��B����y<�UZ[u�����؞���/�������E�MrS��������vY��Ł�i��K#q���w�Td�~�&�,�Y>�\q|�I�o�J!���w�(�QegZ�� W.�����?�G�[�j��P�@�Ku��5�&_|��j���=w�Ǎ(rt�r����a���փM8����X�/Q-�É�Ztߞ=���a}�;��Z���XgB uj�1�u��a~;+]z{x7�,&kXl1���]	<ӧ�*gh�!�fx4�>���̋������U0���5򧰪1�����ѱ�%7��K��{�h�˦7�E�Ђ�>��C�(
����pWl3L#��ke�E*�/���Bc�ə9b�#��"<�*��Ia���d��%�wn�;�'�F	t�K�A^�5AIm�P�M&t\�;��C���Ӿ�����ܣ���ғ��nG��<���}���q\w)H`$|!v\�tCDc����ߟ����P�s5(��ȠB�^��E2��ΞֽS癟�S�$�EH��4v�Aկ6l�,��W�cC�%x����(g��<h�P�ׯa>}?lD�k�
$�8�������4+�}k7�=�0 
e�Y���N9n����{�D��@lM�񘵨2��n��IJ?^go��*}�X����9g̴����f��	H��#ա~��o^> 1EF����o
D�*/v�O1Kl���D'�qB�<�� ܵ9?�b�\9�I�
��_�e�z>�L�|Gu�VeO%�M"+�L������)����dۤ���=w�>%��ר�Ь�.��|^=L��C؀r�x��G�.�5l�JE�Pr�<=3J��[�˂J��\�4�5NdZ���,�&,�| k2�($��Ӹ>�_����3�����X�ZqN@������w�������u��|ƇG�Dd
OrK㲌�0}#G�e�.�t��iY?FS��y6����������A���&}�:�Z��NH��^��Q"�º	�e���z�K؈���8]��֕���le�M�/�^��QBĕ�P�������2p,�����b�Ҷ:�����t*��y����?�\l���i�P[��ࡦVK)�2O���_N�~
�z���#��;�sB[���O>У���]�Ze#����,f�&8����^�
�e���O��x�Lh+5P�٧�����N��X�<(ӫ�8qPK����R)��պ{��[+�v�R�pz����P2�^����_�p�P(�¼1 ��A?�iq��h����X����f|�DP�'v���4괩*�o
�
��q֜�I{G76g�<�I��������ӪV��䵾�(���S�P���,;d�W���,�AӴ�Ԗb�]i�wJ��{>���n`�H�Yl]� ]o�ף�xvnU������j�%f�8jr�&���8h�Z�Yͱ�%�����+C��H1{ݡ �}3�۽TN���U>u�2����V2?��t9xS�a�G䧃����-K��7�r�<�+�(���J�Ss/{�C�
�8im��t_u��E>��l�"f���1��-`m�>"H��!IZ�9���]�}.^X��@*xMx������ΰ�'�n;����7A�g7f�5ǧ�Sѡu�?�T�Ț&��汹���S_l��С	q{�&)���c��^�6ZO�_�&(x�B#8�yb>�G�q�:�4�D�cv>�<����7y9��=lXjB�.���5s�ϱ,*BQj0��p������l����T\�l
��}��(�9�t�s���f���m{ʨ]������u'�'c{t���?&�r�P%����bGy�R��adpQ#�݇6����D,�4��A����L$e���#�dry`@�9�$�Ӫr��N�&ڸ�`h����t�;�Oҁë<%�ɓg�Ǫ�5J�Y��E�bFW��Rh�K�I�e
뜸�����@ -:-�w[2�;ֱ޽�+\	�R��.�X>���D�<���U�WOK&��Ԏ�=>o�.�� ��C"q�l��p�\k�u)FgmwHL`햱RN�ckg-p��BJvB���է����K���\�#�հrh�,>��l��4���P"�1�͠��./�fĤ�Vo�����`�X�M�u��F���h\����+RM˚��C��5־EF��:��� )B)
�i�+6jF�[X���fڧ ���k�^�]�E��]��`�٘��H�*C�c��P�pbVx��^��`�6��7M(w���r]��|Y�݇��ͪP=�Ə��0��Q�F���y�6;��n��zI��.��iV>��^�2�љ����j|��S��P~���\TwUڳ4"B��T��ԢD�E�<}��L�"5�AL6��M_U���sIN=�����1ѥ>��bm���ҡ>H�xE͇ �ph�[� xt�;~~�x:���Ar
|Rq��W��4�Q��kϋ6�|RTwh+o�L�Ν�6݀�P�,h"�H��[�&��y��%�Q�L�-������4�RE8�]�Q^�\GB)���>�&�J��$�n�<�\�$a��SY��������)�g�L����ۨ�xM)�
���$��W�Mv����"�V;K�7���Þ�V�`�|�����7[����� m����!��w��b1J��L�q�b���f���*CY]��?�����"�W�Xf�(�x2=(�m��?+�n|��  h���3��J�ɀw�J�Ojw$5`���� ���!��F?N6�ېA~�K�֨���� м��M�L������s �8cM���