XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���7�p��fc�T��HNp!�͗գ���j0��\o<�R�����,-v��-}�[�^�؀3sǇ��:�H���o�|�V)ֽƇ΍	�QK����z���Ŵ�b�b��'d��P�um�B�rZ�Q�S4�?6���V���[�c�ɬ�\�l���f�&Ɪ����CI�-��6v�v3����u�ɒ�J��:޿n,��~oA�]�bDʇ^�f�PF�~jg��t9�a����(;�R�1�
�W��G����T�!� ��W�.F5����L���$��5�
&��3��:Ŧ�[x����y�&O��K�q�@�:Z�}Bt-U8��'�Vj���YG��Иz�6��^�0%�.	vRG�u��X�Yȴ:{���"�"�!��3�F��-2���t�������bT���[x���E�	�a���!�	�G=�RDF�~�CG�n_~d�%��Q�J?7�:%m#�3	�D@ޥ�
�A���4)HB��d�oF9md���^7N�Gi�ɻ'�Brg���b�V)���S�:�dR�*>�wR��h����0���$�jw��ZCB�7,9������]����$�$����bXöa�y�;/VE�@��7�7��%3��l�d�L@��:�؋���xo�55��5r��"ԹƮ��ɸ�v76ޥ���R�k�c�g�6�@�&�s�dR������^�os6��n�,z����l��C kO�C(�����7��d���m#�υ���p�_��џ�mpT?�XlxVHYEB    5909    1550"���7�-j��^�&"�����H��3���@au-<�{Kr�&�����b���Ψý���c���ß̪����E�o1>�X�T%-
���f Ku�5UR�JRqs�I-*�I��?rz�����"�%�.����솶H�6{+44�ub��k�s�*C|6v��}i?�ʑ��ʛ ��?�>"'~?s�\in)���OKt`����)�����4�r��%�Hރ��6��|�څm�P��yO����Di��a���]�C@�HCE��^̗*������--{�>V�.��K��A�����

w������f�F�!/EM���.ʩcyX�Q���4�)���o�����O5@_�FX�]���b���L���c��y��[��7�K��.�^����� ���X���$�#�I;��"��=�#�����v;yL5[�(�Q���^�
�|4�&��G-dP'����p#�$:�M0p�����+�?̬Z�_���數�O10:b^���Ϙ
`6V����~"K$0��!gj���g=:�X�^�%�v��^�[�J��Ne����-��V� �џ��]�N>��XaT�/��!b)�s�'ÿ����rpwO��I����5�rrQ�9�İ�È�5��3?�
��{m�@ѹ��5�?��d��s�=Ek۾%�p-��A�jf��2�A��7V��b�~�b(/�����yC𺦠�z�H�E4r*��m���8�Lr�l��D�6���o��!��R��X�1"�0��O����5�kk�E���Ha��AS&��B��G�CdAs�ir|h�������_[~O�����f1Dßv	������ �~�	������P�����E�ELL��h������S8�ʤ�n+� ���L��\v�jP_��JހV���4ޕv���?�&Y�/�X~�A��������&�5o#�������?�a8$�Om6�Gx�
��^#�ơ1c�r�*gh�jI��d=S�E����j���҅˦97{�܏B�s���NA�d�|!Zao�"�����0�촓��������MB]M*9{��oN�)�p��a+ ���U q��}�SsB+� �V�5��R����A�3��'VX ��Y[�|�[�@�R�|K�U�ץV�������>U#e/�c���l����݅�V��<�4�Uv��u�����@(U��GI�����|Vqj�N�����	��-75�cU]���$s���y{w>?��V�t8�Ԋ��G�~�b2�2}��]@T*֜�|f���O�1]7��7]�:ʤ���PTO�4��U��5���,�Ͻ����=H3�g-38$!ݒ7�o�[�=�L����aG���I�Ni(j9d �w�3���[q�XD��� 8��*�^��%���������8)(jYYp3�1f&IV:��B�xX*%�����qzL
�����f)��eU駃5�K��\�������4�R4J�B����Q��$اUϬ�XI�>�l�א��"�ko"�rK�m}��[ܭF0f�<���
D��z?���qǥ�[Q�����/�Ə�qw��{�9eB�&w@��
d�)��k7dh9F�>4q���F��o�8�Ȗ>�¤��݇�y���T�l����ą㝞fDK����c��HT�{��[;�ًKh,�䯏V�p�/@�։#�\ q`�ͻ�7�ğ�t����=���[}���-e�0��/��gj`�QS��.�f�z]�I�������0[�Z�Ǝ���؂�B��uP�"�i���,���(?�0���V�۾I~�[�/�u9`Ob4��;��TO��Y\��]���ć�0��\��̻-�Lo����a�)6�/����&y�c�<���&i���oL4���*�B
�;<<�*�+�J@JmO-��0:s&u`�qG�ֺq��x��ys��+�:���wmWf�<�ު�8��n�Ղo\����iHA.�J�qL�V�Qh�߳J4*U._9X�N�8i�7WM��rk��`p�)Jl��jC� ~���t�闪�6Z�A�����m�;�vM���<����=���n����Mr�p
[�7�BJ���
�I��m�V�r�Ox�C i��D�"u z�&!�i�W*]c�6�.��8�|ɄŔ��?��[�f<���#K,���V����7l�e�I}!�ѫ�6�̾�_c�����>�9���@�s��nf�f�gYc�!���,5 l&��LR��(7�9N`�H
a�]Y�����i��00����q�(O{��ÿ���c|���q�#��Z|LO>]<_-B��R�R.P@�tɜ�=�~�[�RJua���B����I^#@s���H���?���o�	(���m��p��.��qf	O8h�,�t>���V�f	
�z�����qs*z�M��(�W�4�p
���$�Q'���7^аx0�A[����o�Yd�!?���/�A��ߎT�Vjx^MS>�J��ߐ �yT+ ̉$or����DtM��m~�u!�A�Ղ�ui�ڴK���z`��pwθK6��C	��a~t"�8�ޠ�ԭ���T�Z�kQ�!m"�=���~��m��`�j}��E����� `�>�?-:*>�l~����mX U�p"��up���$+}v��qS��1�A��bE�I��'ƛ�ω!�i���f�#�x�F�%l*�cs����H �➻��b_W�Y���|�����l4ٓ�a��B�7�<-��������:���#�Q��o�_��`aI��p2� ɛo��H� �1Y�V&�'+m`�M0z2�3�
���D
Q���I7U���<���2��\�>�-�ᾤ�g��"���9�~Ƽt`�.ֶ���Ɠʟ@"���5/Q�����{$���p*۱���G]�����o�`���2���%r��v��Y X�b�s�oE;4�PE��%?ւ�Ig��q�F�$+p��9S�]����Zetz�v�F�XƷ�ߏj
�6Ƌr�����Ç��ݸ �E�{�
�ѝav�4�t�l�	���s�H:���Pt�g�Yn%�=�+}��&%��e��&j��yXH�aԋ�[����\������%��a�����������o_PQ�����Y;\�A5l���D���BvM�`bA\ӦET�1%|�C�9Qш\��rF�sW�r����aH^a���:e���d3e��T'Ւ׋')�g�r�缒k�� I��}���S�@��ܗ.^�*ۓ��I�?(��:a�<����_.��
+�5k®uT����#�q���u�����'���!pk_Қ�r���Y@[��e��s�����% 2�Ƴ3v�zWfY�,�	D���6�c��x?�+Z ��q�ID�$�py�9IAD�4��L�����p��u��lHȻ�wf?�͉�}wTT��>��g5�]�n�y�@gڬ�S���&)1@�"��_�gʐ@��p��jI��g�˾�np y��.x������u��q�Y8]Zǂ-쫴�:0-b~jzQSRY��l��X0������;SZ�3���T�ƺ�jy�*��L��F��������P�cd7�,�oZ���ֈ���
��i	s�[�e��V9i�Y�6påj{�	Z���b���+��gHAGLXZ�"�e>L^�����������g��^��P^�f�Ie�������'hX70(��r��Ǿ�=�6["t(a�GsR�o����?~��
��cC�[����u!�""S��b6O��$�#E�ѓ������p�2ڏ����2a�e���� ���0����s���2�\i��ȶ������w�1��n����ժx �X8A$GR��:���yγ6퍴Q�%]��%��H�J�D��Ʌj�g�j�Sg��t)]!���<ԋj�SF��G��:�0ؕ��ru�4` �"��.��׍��N������ysU{�k�k,�[����a�a=�z�ȓНN7_����U��!hB�'���F�9w)q�p"zq��׏Y%��azQPx�s�W˼�N����kIYh��.̸)(
>�V�Ĉg����vA�̥�q�\ �d��s�B���h/b)ߎ�	��mv����K^==���S�'�=ޯ�QZ�+�,��I��������N�	��1���$x�euR<��8�N��u]>C_,�1zC�'ֹ���Tx)�nr��i�`K���}��He�в�TQI������Kȸ��(m��S�VC��[Ju��-�9/6���߹4���i�xBs���j1(ii�s��'���PN�=S����ܤ��JZ�{!�X�RL��	��{�Z��� *>`����ߎ�:lq&=��Z��V=TR��ap���}���g�k��3�O>� ?b�;�9cCj�9�������c��h5d�/Z45\��'��a�xPL�M��T�;��Xs�g� $�D�P�j[��QhW��uc8�D��𠼫�p��= �Ǽ�G9�c�`��RҚ���H��{��-����xh�E۷\R�E��rH�K�m��[;�q��3�x�`��ߗ�/g���L�w�T��"���f^��闦�7B�LQ���*5�~��2��8�Ѐ:�������f����{+{��@���FR��$Ċ!�<p��%��m��%.DSʮI��S�!O!�k9�e�q4�1:~<�Y�&��������[j�8�#��
 Gw���~�)��C�3����8�k� d�����,�/f�+ٷ��N�O�oU�d�+Ħw�0r	��B��>�2ʾ��Ɉ�����lr9����t4	����d��݅Q����=Ϩ-�猕\q5jJ�:G�1iV��y0%�g	bZ��mK��[/s�V� Bd�X�!��Z�X�XH�!��0��u�b���`�pZ�`��`����]^���
����)�&�U��vm�����h46�jMv��ݷ�f�XOD�����8Q�=�u���@\�c{�� ��\<����K����xD�g5��e�hmVk��X�8�+͹9�C�\QY�`����E��,&���T�s��RN��^�ét�>/A�_���~���+�9���G���� �K��A6��u}����Ƴ���} �0�� g3Ӂ@��#�<? kW����{�e��EMd��~&I3�&�`�y������8��b�>#EL��� )�7Y���Љ���Q��Z��^���XyH�]7g��0�W���o���Fg�4$��pt|w:���n��|��a����΀m��~e"���D�۰!% �_�?��i\����H��j	0ļ�@@��+/�bf�=y�7�~��hR�t��^��C�ߩI ��]�Wl;�&��ò���m�OQvG{��Ţ