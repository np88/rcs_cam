XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����B{��Fzc=N��rK1�&��|zCS������������Ŭ;=,�,��c��f;�aJm�J��\*G4�����muD��ca_?9��:)����V�Q`�L]F��Bw�bZ�a�&Aǘn�[-`T�LBz�.J��s��w؀�F.���Bb�}��#�[Χ�r�K��P�G���`�R������q��fy���B˅�m�Z�!�n6�J�<Eή6��(5��(�СDPH���߉\D�㋖�Ό��-S����^͍(('�|�3$ӡ\�|@�M��?p^t��U��-���[��O�斛~��|�U0��헪uMyw��иRݘ�h9Wn'���ʲ:�R)��̦2�O�al��m��amQ�D'G|�S�n�g�ـv����D�W�$l���|;��[֎�&)�[���>ʺ�X!�s�e(���91@"8Qҙ�P�.�GX�BA�$���_ՎL��L�̚�)�˵z��1�h�M�P$�/���g���S�l�w,i����q
��� Q���*�7��y�V����U�0>�F��4��+ ܡ4����yKQ�Qz�w���gɜ�r����W=�r����~/A���L�ɢ��ъ�wL�}���7@ �h	�#�`�E p���d�A©��g����-��t߻�乀�x�����$�eLcx�eOlcwx�q��|�b=	A��i�lo�@���fiJ�r
��?�����k$3�Asi ���0�&o�H�+?��iQ{�K��key����
�:y�z�~�XlxVHYEB    5694    1280U�ğ�*%M&�Ҡ���飠��'��Z	?�0l��T6*��N�R�獵��q(1>�k�͌9%�
�P�X%�i�{9D��?�����2v�bj�a�&���d��E*:��5�iy��L��i����9��<�lf���R�-e��\/�?l%���ga�=4}e���_h�{�En���J2C�;R+i,�
f���G��$"tGR=|�+v�,(�#=r�Li��c��ʣ�]7�o��a�i��Iʳ�2�y]�;w�X;e_�c��j_��"~��DCQ2��x���du���ԕ4Ӏ����	�h�?�՜ c}�)�Z�Pʭ��ˀ��F0'��=�9ìj @��C���M�qV��Q/<6���0�{��b?�9�@�D��Sɖ��!����|dS�2��������m9~��*��;��
.����f�Co6��䭃K�DH'j`����S���j�h[�<m��TTh��bIϔ����4}��?e����@��%���D:Ӣ���� ۈ�y �����寢�p��Zt>b��yVa8���=�K�9��n�� ��;z(�r䍤������-г��X*3&F�ێv�&Mz��{�_8�D����k�����zE�DT�SKY�!MI ��JV��M�a���:TC�h�I��@��S����9�>"���M�]��v�8���v�����r
iJ��t�
��#���_�8/'BoD�:��ˋ'�j6s��/<	>q#�$1���M�gŒ�@j��A�>[q���<z��@����*1�
(ֹ{�������oO7���?:y��I0�iz��D&Y%j�l�SaC� ��LOfQ�o�F��|�iw�����.�j�A@E����j�kI��	����W�ҭ��B�J%�;kD�]��6k�	����U������ ���($�/�g|-���
�G�8@�d�ڊ�Jђ��S���3Ӣ��X$	�ܡ�Ϻ+c�eK(�R)��=����d����Τ;���2�Q�޸��G�W���JܯO��?L�`H?�l���a���W�[�pj����=��$�}ܖ�>MX�ꘇR�M[oU�����R�/��&F�s��}NO�6��w��G��(_�a��L���ͭy�r|1'r�D�[,Iq�/J8=cy�Z� �� ���ꛬ
�*^Д�L�S�z��3�S��^��)7�W���X>����B���T��G%qL���2���ho�i�S�� ���1�$����g��أ�[n�o�J`��<��ԯh��o�L.���7LY��@q�l�:8?�3?ˢ�& ��;R,#�z]�pv]Is`��L5�Q�i,�ë8� }�#s��/�i����+Ct�X=���я��w5zя��>TW7�9s��C�
��I?n���/.]CWX;~{Au����;��Ĭ����u�[z�&]�V�EäV ���)ˀ�V�bKm�a�`y���E����o���O�n�N
a�<r9���c�L3O��fJ7�4*~�$��'�v8>t]Ї_! ��x�.� C������j��5� �F}b� ����`{����y�ж�����"��j-@�$�vo�׸[mb��K�@�DgE 7��S�
�eZ�k	Ia�ڟ��AR݇�#쟜�W������Sbͨߕ���X%u�����"A!Y�g���Y>.���[8.9��D	p�?��2�ڵ�7;�y	��Q����s?9t8@�J�╚�Z�ԋ��7e"��0�䢶�kZ���>���L���`a-�őt�)f���(�O�E��dgbo{族#���FK�'�3�5>�;�l�=�t�'aG��:އ�L������� /-�%Iz��J�e~O�v	n���1��'E�Q�W3�,Ern>[˷�;zU�Z��UHCW"�M���޲�	���66�lյ����r���c>�ڭ��Z�n&�{�")��5z��a�e�5X�ݯ��������VAD�%p��~?��n�<X�j3S����jW�v��?�=���Mѯ�o}��sͪdI!�qe���;��*W�����N�9:F@v�v�U��z�������҇?�Z��8��)�E5����ٕP��f�t�ů��|8�Y��c1�J���A�Y���_mɢ�H�f�ľ#Z�iJ����y��b��G�}zj����vg����`yo�� �݅}�-�����[��eV��K��C��}0��og.(�[)%��y	�zv��&�?�9��P�d2�����<h@�d7c,.񆴅� x���wk�g���?��P������ђM4��V�P|�'��1ظp��g_1��)Og`&E^�:|�:ߋu���b	a�c�+����0(�%4��ű�hq"w@�� �WXh�~T�3�5 ����N(�X9�{y���}Ϧ+Q��Y6��t�0[ �6�;�<?�u&�׶g��3��+_ lb�f�����2�r�/X�d_�ШI�FK
ZD���Ο���L_n������! M�lCD�5�:�W��/w�)��� ?������R=
�N	�,l:$��b��x�����"�����^^�g���?I�-|
jŬ.�F#?��A�r�~i���L�9l�A�~�~n>W�A��Ge����E��B�J")ځ2N��J���Z���_����_�b�{�$�d⊙�����%x�x	H�X�CƅrX]+�<���nU�N=.Z��H�,���av�s��cEI?��£�>2��X(�@�0����>}��W�O[U%m�Wź�6��cV�l�?+��!t�sY�:�&���|0�W�|,[�Jdb�L�����?������04O�t���6i<��.�0'�r�.d)0w���-e�(V�>`y�Ү�vKX���ع����a��חͪapwJp-�3X�A�Plj��m�K��ǉ�1��I�3�P�;w.0ѭ��me������DM7���3c�fL�a�������6v{�w[�����#3��wt� ?.E4�n�wٲ�ۗ�󴜅���v�Ғ���_�S>�G��+7�i$�[�ǝܟ�b��ӽ$�Y�7^뚳�M�u梘¶�L�3�3k�x�n��A4��tw��ܼ�8i�8�&2!���qx1�Fվx3�-�P�a�z���nC�@���.�}����]7��&�S����v�������b�3!�n	Ov��zh��9�?^��:��R��aV��QC���!1��p�<Zf��� F��x-W}�� e�?�/��p=���kb� ������2�\ ̰5�3�@|��G��It���zD�#=}�4��kҪ0]�̄���u��>C�r�*V�v"=x����]��Í�� ��Eȥ�`�s�5W�P�*���fZ�aw.pm��a����ǉ�P^6%n�|]~��&#�~�Ư��`�G�YA~�ϸ���^��d������=Ϩ���K%V�y�!��vs#�AL����h��PFC.H���� ܟ�$W�v"�����	54:V5y�ݍf/�)�ޏi��nV[�=�`/��槅��aF�п�7��1����6�(����"i?qe�T�l�j���׎��0h���<#s ��mJ.�GG�k����$�B���/�#x$�(��S)�@��I�0�_�#���/6��g���Y7�'-�Z��6�٢_&�:e�DX�3o����VV�"�Z�V�6�_��=�oV��W�����L@��z������p��	�鼼^mè>�ŧ8����[�h�)�X������4�����}���[j�#�&�`����nD$�9�;���IC����z��#��'����>k�mFp� (��<�A�ǲ#ȳ�O��g�9�D+)������􋯆�_����ڕ��=B��ʶNϭ��φ#�N>���E��{� ��힄g��qF�, O�?��PB�L��W����凼P���-�.t���\�.�"P30�"�l���=�(������N�[A'SaU%���iBK�V���u�\�$@P���A%��Q;�TJD�$n��Tt�hl �{I�S�ac
^�E6H  kkY�{|�eH��"}��� Y���&�����gIHQ=}$���Z,���6�{a��az�����:���)��TuiK�O�r��~������w�P�uozr���3g��6���R[wCe����X��l���H�N��[y&��}ɉ�C��g�5a�ecQ���m��0�
�y�L��xvdr��v�������Q�+\Cz	�3������%.���7i�\t��Z�$�u)�Δz�¶� ȁ&���{��{����q�E�I+|W-���Z<[^��4��^N��Ry��=��D�(�R��;�J�{ L3��ú� �qn1�c@hV�����I�8"8��c��"�<���������n��>�VՙB����/訔K~o|e ���lV}�UM!������vW��û�Qۤo���#�e�8�����*�`夬���ތ����m�%����ϔ�U3���1�\��qX9��n"���>у��T�2dU������2����)��5�|�
J)Z�c�"���#�F���*͝�.^�d�\�S�vd�fـ�XX�����T�a�}��r