XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���ة��D���u�ҝ��+��R��G"ؾ3�⸁��m�AŚk��4y�0I܅p����o�gV-
,`Ϫ
���$eI^癣p�1�|V�j�}D9�����l/��n�X�WY`e�è\�;�*#�Ƃq�m�C�,N����=�"�E M�6[6i��u��i �'!Ƒ���EP�����J�e��{8v�L%?�O��R����#���pN�z}�z)������/,�^��!�#ry�ėS��\4�oH3ؐ��|����n�9T��RB^�XBP�����d���'�F�Vtt�F{as.���Q�X��6 ���]�k<K��9�K|.�6s��6M��}�����a���7l\��5�ΊЈ���ꂈ��td���H,���
�)���r�~� ���_q�����)YzK���8����=���.�����h�����	�% �*�����Fd 5P,�O�J�s�b��?H6�{+��m��L׊3�R)��KJ���G���W�?�D�� =fPc�O�����c��Ғ{���Ό�(m~�>_i�=Rh�ӔVi\~R1�1VY<�]}�t:��^d��L�!���&�4p��  ra)�Οh��)*.U	��2`�VyB[x�<�=�䞪�}ܕhi'Z���77F�M��ز��R�e� ��ΏC��i��rX`C��LsT&+��g��#Cau��(`����0�p�S�*�K���73u����p��[ޣ(P��0����?�XlxVHYEB    fa00    1f70W2�q1��W�T|-�k�׺\�� %!�MᵟJ���~T�����d7Da�ztj^����r���T��mN?igXc):��Oy�g��f��Vʍ�k���,re?�Z?�����!�;ߌn�Xq@ӯ���@N���k�7
�o/@[n4��Q�R�L;�n(�R7sD�<L��3��:FY�+����@������a�e�F���� ՛b#I�j$,�����"�[������Lˠ�9y�BS�1aEy�ͱ1��nF�8
����a���pnvS�;ͽ�E9��A�]R# � n����!
J&�YE��x[ղ�?�L��o��9fu��!�6���c&Y)JT�ۄ�,_[[�N�W9V?F���֡�I�MS,��e9}'&,j�Z�]3��,���ʌ�����e���L|���n��A�D�#���!暼Y���i،��������`�ա�ɟ4����?0����B��+s5������f�˲���=�풸�ΘE�s����29����K#eRۋ�tV��A4�>d}P�8u��>�%4�iB�����ؠBMgln�>�pn�:����!r�[�<��Wy�'��係�B��f�����
�=)�<�Z1+�q�BҲ/Z	e�PeԈi��������rjk��%M�3$���--)�_��3��v2G%���� F���q�k܏��f:���k���R� ǽJQ�mz�|̎���2�w���P@[=�9j�+� �wo?�.�j
mG�����Ԇ���C�Y�#T�Y܅���9@�T���h���L�_��)C���/͒r���J���609ٖI��r�#+��fs_��+�H���M �?#raA�Ql��!���(��P\�
�n8�;N���R��*G;�R�WY X�!�8b���/N�K�@��� ���Aw�-;�T�\>��a`�I�32٫��_k��I��Bg��/�̊�D�TCx	2�:����w5��Sq��	g�	J�ê��I����-�3��N�C����q.lس8`*��H��K��j�`w8��Z̽��E���	����Z�2�����7f���18Q�5YD����.N��8I��d$������)�-LC�HqZ5|�}��M��� S��hX��Ċ��(4�ǂ����#�p�?ldTY�Ξ]�[|PD�h��x��j���C��F��,����A��z.��a�3�]k����j!����#w����u����r�]4�����+ViP�\����S�&U�7�J���^ƻ�j�	v6�����O����%1�Z�����n�
i��j.���*�uB׼.	*�V�_?S;�,�.��K�&;�s����?�:�bS�
�?e�QOO�{чϱ3�2��&�ҳh8c�h�"[�M�m7�f�߹C] �E�nX&Bz	�9�6�O#��i��÷�,!U~�.�J�jƎ�.�_TKY7F~��"�GO[l��=۶3D�R=-I�n�[�|)�]�9����y�������?���u�9y�ݪCLja�ۖ�i[ȱ+軦
&x;�Ȯ=;M�}]����
�!F.�����ʩ�l�#� ��k�� �d��\6�AH��}�X�����״Lr��h�(;s2����;Tϋ_ޠ�׆�Zz�R�U1�gv!�m�ab5.��-�҈�%H6�Y�5�P0�LѸ܆�Iw��a��;�9w��pG�#��P�Ee�9����'��q��EF�O�YKe"��J�=)��]T$/���~�w��I�W�Ī�Ɵ$P4E�B"���W��`���N�-7T�~>��T�+���<�xO�	i�@6R��Ҕ�ɑ�M�w��>^Q��܌��˻����`�4�)�
٪�pc����T%Fáh�����%�$�!���ҩt� �S�/V��t��ށ!d�vP���4$B`IFtQm���9��b�8#k..=%����O�0��x��b����I�bt�E�����WU݇��VA듘rRPX���ZI��0��3%�9G���Ԧ�����4=e�1�wTM�~t\��'�ҋ��y��?ӷ۱aL�9�Iu2�B<jVQ9��Z.`��uv�+��@Zj�ؾ���$	F���@���+�a8�{@]���K�����1�x�1&(���PS����!pY��X�i]à%��L��!G�v!�.o<Bת,r뛿����:g长�j/�$�,�\�F�h�*@I���8:3� 8`�F�����D�v@N�Ъ��nn
��0b1Ɨf����v�@�
�d��d��fr��-����o�w = ��qАt�p����&��Q�)9.��I�o"KE���=ٶ��}��;P��.+��Ţ��ڦf�7|j�J}6�r���@�k0��T�Zaih RX:�
���A�@l��W�j(~�x��bq��Jo���WP�K�ܙ��u�e�A6�7���'� ��w4�t�@�3I���Q�4�+X~�
M��x��y1jp*��W��f������-����.~.x�o=�
0u�!�����(|�	fA�rJߩz,��&�@v��V�ȼwSП�����^���$�V�Pyn���R���Jƙ�,3��Fx��ѵ��g���Q^ ���/�#i��|U�2��:�rCm@;6
�E|��8H�˷�n�D/�}��(�{�G��"�^��R"��7�
[�ˈ:��^F�
�ʄRmm�u��f�L���'q�./�%=�IS��5���w�ѓ�`�G�0Z,3��&Ǳ@�+�Gr����j"�I\�߄_�5�v6��Ŏ����L OÀ�����_��\B�M���=�&�OlNg�-��xD.�rä��s�4�SR#�ۺ��Hu�]�B=�|PJ�Jx*�F�(��րs�U	�ӈ;�Ӊ�8
|;K���OKI �OgD�Y�5�R��7Y�9
�ϭ^C�A��^�8k"�'2=bY)1R��Ί���-��+=d�{>B��\��������tuNmq��TG��P�
!m��Q�`&&"�k. =Xn"1O�a~(Hͻ!o���z�4|�h}|�3����<�k�)�l�юz�T�<�6���B�DΧ��1<<W��',T��Gz(<��؆:�>��2���Zc�U�%��}J���v8��Œ���K�;[F������Ul�"�4��T�V�Ax���l�#=+����U�~��!� �H���˙`/�[V����܍I����G�#G.g��?45:^d*/��rk��y�d�r���n����B�?��C�����X��z�DqSv��~
�
'�h�ET\��C\I����y��;u}uG��2�u#����30v�j��φ�U1V��l�X*`@��+���B[�M�g@���`.���Ӛ?Q���Ӹ0�2� �g�@���"�0�O���*e���˻#�E5��5���u��FJ'ݴ�Y1�W�s�9BM����m��[m��+$_��}��h!���Ao��H����9�_�!㪨��ɝ�ǝ���YT$���
�?�h
�y��H��"�����e���TVl~�"�i5��O?5[߅�[b�}`��"��?x����
�F�ܣQ�.l�!"���M[a+5��HQ�˙��-�0�E�[G]}b{N��E���/u��>i`��_��fs��N��m��z��� ����o��q��֢Ks�����B���)=)�8⨨�t��7o��%X�I[1ΈG|מ�4K����̓
?VH�(���ºA���*P�f�
Y�xPl�\���,�
�2�GP��䡰��eQ'�P=!п7���}���,��Ķ��]#�R<Ј�J=U1Tݧ����2W���:	�

��Ւډ��L�W l��T�,|��(<��ݚ��2c"{��>MW�i��T6�|�Ne��>Ms/�^`	��T�7��- e�o9��Fi�oE�%@�(uW��?v `�"0�g�R�jq�OrO��E��f�U�Q��*�O%q�'��V�W&�Y	.����X��^s����#	Mq���4�Ch��)���ve��6'mĬ�j��-���\���$��pT`��}����%~0s �T�o��g�X<T':�Ф�>ʤ7$��جO.����Ξ�7q���<;I]�/�|ܠ»O�'�4μtt�A�5Pql�vxk��J�E�ə>���u�[1fQ�?��9++��n����<�7��*9�[[��5�t2�	�q^�`�L �Lz����m|��סmb.��n�͋����ۍY<��?�,��3�Vs��]�wJC7����8�,�c�4]k�˳c��!�g!�0� �nギ�u�T얻TU3�"������Gչ��G,�!20�{d�{~����&N|�b����~I(���W�{�� �%y���ii�c�$x{�@$6� ��"3a�l�8��#���*��*Ĕ�la�Ď@h�|�!׫�-�yr�Էvb��a�?����XO���W�<jƽ��9��²`�����x#��L�K]��7�����]N�j��ً�T3�����%�WxD�+��W�a\�4ZH3�^�-�2P�{v� 3:��HNq�V4�'�m�N���ѳ瑠4�We�C� ,�im���D����-!�Dy�Vq���Z1���ϯœtyH����"ks^2������"��>݄��\I���>�N[�ņVF���4�bW��>,ۺ%�u13��������B�D����r�ޢG��������	Yp����ObT��Vo�%������{t{���c����͚#m623΁]��&/ZG�Ec=�g����	�,�8�Ԭ���2P���|�N��:��1�G��!�{8�l`��n_��arw*k��P�1Ȍbs�y�[������&n��㻧�}Cg����A�e���ˁK��X�[��W{����w ���,1�b9ubx��u�\����a�w-_�>�@�Ð|�"�G�3`i8��ؒ����	��(G�F,�R\�0����,������rU���)�h{�������r��B���"�����̓0�����PA=�X���:ތ0}c�S��g<�c~�H5���bY�U\��%�%a%��QX��!��m��T�l7���G^���6ɂE��)�5Ty��ӷ�hQ6�60)�kR���'��$��+na�F�3Y�d���'�K§�������c���+��|��#H�W�w�i��<��(�CР�%�@\��,!֠;��������}�y�`� HW���%	v��G�W�n�����l�Gh
/`�5t�Ͻ{,1=Ͷ����l�mHo��*p��⯠kțRQ�ץ
;G��j�f��}��%�^�����S{�W��"M.��b�W �k��wԃ}(ƞ<�}Vc��(E^Y�k6ę(����0�yZL���T���:'X���9}�U�yk�z��}�8# 2=/��O��}��w��t�bwo�C��&D�(̱N{����c�޴~��9I�9�6��M\ L>���,�p�{C�"1��u�c��|{�\���q'nM%�v�K�gPMh���=�ƶi~�}����`td�n]O�-B��)�#��M�L�g4�'�_l%M�3Ŗ��Ox���{�N<�,
K<�[�F=��E��TIrqL�*���P_��#�%�^ǐ좼�c{���ᘓI�7М;$EE��|GT��?<�wiy�n\'����+�w�Qя3�{���z��4���ZVs�J�5�~M�Z̗x�! �/j=u2Q~<�q�xF�&�Q��bΥo��C���
��@v`���a�*�����]��ɴ�7Z�3k��L�<��j��r�99��n��l_�T���(�&�Y3#����/e��$o��"�d	-�27�w{iMsUa�m������d,aᎧ��M�R�j�����a�ʙ���\v�=�+4��$�t���zB�
>��di�pq�̾���q dq�^�3��S[f�r?y��\(Tu��V���P�Y�3�j��BK��(B�`d=/]�1Kga���[��3!��c���3.<�m���q*�^��c�%_�A{Z5nS���Z�
vIcT̒��:d�+&m����䀯;�-rĿ=�z>sz!V؀C@��!�^��{=��`+/2=3�-��E�p�]DE�>��T�C�X1& `g� ���q���U���oRlD����n��e7$"@��Ć���LES����h"��M�%Y`��]���{�;A|�F��bumٱGП��yD�H�~@�}M2�'���rM#j*{�I�W<���Z$s�p��)������:��06=�Qf�3�2��E�GA1�� ���@n	@$H�	^S%}Tf��y���C�z��ճ�:����<I��j��XAj���ԗԘJ�2�>pa�05]��1��������A�LUc,΄�bw��B�y!���b+�<�����)��b���׺9��9��.�)������FF��sO�6C���aOteT)kG���z��{30��q����_��'p��������Wk�+|�s����@�މ�">�ڤr�@Δ(�a�r6c�<oij�Rb>�� �c�L�|�E�$hc�s�@����{�~a�\���]���do#�ѫ��u�"	�e����xls��vџ�:2�H_D߁�;��_=
\��io�ث�K�G��e�%%d�tEW�S�b��J��N�� �ԘW5�K8|�]@�6D�f��G� {�q���ĸU��q~�ɝ��zf���B������ǻQ�FC��u�,�M�鞕g0�y��{ƽ�"5Ըƚ#�8�����+-5z�7���f)X���e&}�̾:��fU"�1����!x� ���s[*=�8�������yMU�ж��ͥ^�t^�5��s�Bz�d �|�Q�wSzl���.�V$3��D�T�|g1�;\A�d��%[Ѿ���fNڼ��<��aKޮ|."�Z4l��ر������'�9w#��������G��u��k�{F������L���d_3#������|������w�U�?��*{hk��N���\��=|�l�)�Ĳ�)_��W5>���>4%t�h�>n�7�'5���I|'��x�w�H�:�E��)���m>�0W)e�=EW���~V\��C��nΧ�	���L]s�ˁ7��` s�y��R�+�x���n��D��zR�h(]��lL'L�d�Ղ�K�q(�+�ޮ�&�wv��5��^���23�SC�A�awt询A��-������3K�gEK���\��$"1H���WB��1~�3�)����r#����D�YzIӒu�x���X���� e"jA��.-6��eN~2�Y�����~�J���1z,-I@�쬅�}C�2}�-lI	�{q�ඍ<[lXƕ��$'�*����mW��ñ}V`=�Ǽ�G���'q���tm�a���X%yo[����4^Aۘ��NF1)��E�Fo��N5t�Y?��5���»ԕt�.����hq(�|Qy�b3��Z��M͙Wߊ�N� R�cn R}������@������HֲIh�%�6�eNF,DaOf!P*C�Hw,(���T/n��d~��js)ìԍ���!00)j�g]��s�?����
��H�4����Xk��Z�e�])7Iq��Al���}�P�Y!�-A=��Ŕ$�&"ܻ���y�e�F3��R�b�6m����SSv�o���cRpnTF�lt# ��	Y�6�Oq�����;��c���MY�C@�����E�9Td���H��&+iM7Iӣ�Fg�t��Y~���QV7�}S@��x1 ��<��-�S[,AKڞ�� Ht�#*�k��,l����w�PS�dјSm��j<nKO��r�:�XlxVHYEB    fa00    10c0;��g�f"zj�:2:7�<��wrDy���}LxUq��%���ȭ�bO^�:�@6�4����,��� d׈��]���W��d��`xF/�}+��0�0���yGKY\;.�Sx�/L��S�7ނe�����K$� �kZ�|�0�g�-�{o��W�״ _��H�A�N�Y��Q��1yx��[�����%��M4r
��Z�����I��]�]%�H0�M�S~��'K2��ե1���#T�5Q��j�?�����sH�4ÈX��;��4cPqல���T��&u�.I`}bP��}�jrC>p�!&0��F`"*;��ܴ�7�|��%iމmX+ی�þR��5�'�2VW>�����\�WI��R�05,�u�oC:�gO;^�☷4vr��U�cŶ8��Y�=*j���%1��dA0:�#�i��yK���4��E̴B��m�H���Kz*�#�
�iI�O�J�6�j���4>���A�+]}�ۓ��� ^[���/�"P'ʔ�ow�$��^�g6�a�@�Mm͙#� {���Q��)���v�h-I�QJʵ%7�ﮣQ_�,`$JL���ja� o=��;@p��"t��~xC�W&�|�ͷ�-j2ԩb� ��v��kGM�g�oS���c���\���t������1��(CR�2fk5������IQg�<�i9Љ��!���Z�6_�Y�(�M}0��Ru��Q�|./_�3&��j��0��ȗz*������l�e����J�3L��.�΀��AJCĿ�L�����G�!��K�öNҏs�8�ldy�2#��
4�r� |C\�1��W�tA�P��i&d�;.!���=,�>�	rͣ�z@��yƙ3����Ԇ8ʐg�����~��%l��L$%hCnx�O����a�+z��H�3A|'m�
��ILh�c�}�DX![ �25�r���d�,���v�������X���nP��{hU����i���8s���OCm���������o`N:A�۹`0fQ.���^���V&�Lt���A�Q��ި�!�/�jh-��W�Eh��C����1Ş�4On�L�Z鍼�F�W���{v5Zq8F!ґ[���1w�L�|*�d���6򿑹I}�B��h�l�}l���Yb�Co����$��V���ܘ�-gs�P�븕�.Xo��/�%ېV���|���(�ɛ�f�8�+K�GG �Q�ћ.���p~�S�`˖�h��-9�Ro\� 4�����������ΡM!.�d�P^c�NJ���}*������;����F��uiuI�Nk�Vhqp�uǆW�M(��q��7�`����x��N���]�IH���t?b���ix��@�����.�SKS��v˙�쉴�D�%<����Z �}(b�V���S�^���WbqDE�.ܗ��!�Bf��<�Rz	������kO��c
�7��� �%�xV9;J۫S��x�b6�'<z�g�?o������~�Q���o�s	���W��Ww���J;d�IE�M������ HC~���Z^G9��rS���AuϾv���/�K���E��1�r����oq�Jc����t�d���mCf��3���<}ˇ���	[^��E�j���euC�[�Y�_sLt$$��4�L�Z|��bXq4V�\����I� [I�z���p�lya� dz��(�����Âꃭ�u���y��f�T֜Xj�ޚY/�qK`���"uu�f��SX 3����B�C�*++IVx��p|��G���
u7Z�Ͱ�N�ܓ��_.��^YT�Ȫ�Z�����d^oo����V��2��2�h;z�ʚ<���Gv�9Ӫ��nˡ��*m˵�hw&z�ȼ����d�=p���޼�E�g�2���.��-b�Y���Lk��sIKw����9a`Z��y�_�$>k5 ���6������ڽ NR�U;p�����2�t$F8�g(�I��dO�g�8����~l�Wq8qi8/�X���/�2`�MV�Ҷl�;;�M[�����=����ψ%���WQ�K^Fƽ���Z���/����^k����OdM����t��ѕP�_)�/\tG�2�5��<�F�0���ƝW}�'� ��4�RN���:���<���ku�ts��
Q�j��^:�H����8"��{"��,H?x��7FH�������0��(B������Vy����V��3�^|���j�ʤR��
��}?vb8�#�J�6�I:��\
�Ww�y/CM�s/�S40�B��Sb'[%�����t%!Ny0�'ړ��*v����CH��~��9�yj<���0�<:�
��]�˖*�(b��M6�t	
�AS:��	����೶��z}6�x�p�vDID�a"{�cV�Q�@�e�g���g�L�߈C�f�6�h�O��b�~�ͻ�2���D�1n8q�ն�Z�h]|�ݖl��!1��n�v�(����Xٝõ"r=xT��x�4H�����}�	n���d��:?�Y��U&	�C���Z��JX����ß�ߛ	įeU�Ȁ�����d \�����R��"n���T_��i㒛w�*E!ɻ�9�.��v�Ybop��v�ߵk:��ݧ���'zM)3{.7���>���&���A��>W 
��^�����^�i�J�W��o�Xt g�G���DQd*�@⃌��w��^*�����5��Ŋ�ë@�������u�_j,rm>���O����aT)�K��'{B��e�@Okq���؎�:�q:e�[9a�9Ѣ+�xӾ8��qFq9\q�XXΈj����<�����ihvı�ٗ]��M�m��`b�t�
V'��fy�E�����z>�hU�?��fX�l��H�V��j/QV��4s|pi�O 촙��/C!���g��Ȣ<�V�ݕ�{X���\b=Ɏ)�m��K܆�#�\ǝР1�O��ײ��җ�)2�3=j��9��:�k��0�}�-�?m3�N
�}�%�,�o�Me��Oe����Dë�y�~#� ��'��:�_����.9��pk�!�m��_�n͝uyx��NY׽�����W���m^�K���S�:����fPb�,���"��>���.5A�%�DL�v
�dm]=�9�w�qcg���"�(���f�e�mtҍ�'rY�m$��Z�aK��^�����Az��k�M�����W�꺊74�aU,j٤-b�(8�u*�@�UC���P��ИM�O�����v쫌n'�L�{�"�H�����KT*]-��0=\L�!���\9�.�bs��6�4��O�W]�^b��5��%���8� 	�d� RMk�N���o͝3��Y�:ƹ�|���� bM��E��[>V��������W�)�;�9�	N;ob4=���Oe�P�����H���)��ė+D)hIL���C�]0y�����sG�C῰Ȇ-��}	�E�"�G�l���ܭ�^7�U�4�'��r�'�{7JI��p܅��Q#,D��M��T���;�Y�%�[��/�Цu�ֶY�*9�ki���V~D�U��������	���@��-wv����z;�:�⒞��q.y�S(@�(*�����?�-r���k��o��j�ǋ����Ȃ׫�P�����K��%!�<Z�M�u�����P�W�.M�4���K3�t��D��p�C��s�DkDܬ膐�"����c�UN�B�g��M�h!��YmvYy��>���*/q_*���K��֋̵�MpZ����pTf��!�d è��T^��kJ�O*q%3�Z`o}�5����/e�Y�&�������6����#�7k�9��|��)K���'��{�0��DX�d/qz5[qv_��>���TO�;�\wZ��v�g#����� |�f���tԠ�Ql�H��xL�
^.	��S��oB/�2��+�u�r{�r��%&�0N�ZZKiM���''Y/�=a[�к�{*�q����FB������<߾�۵l�r�lw��/�_t���~Z,\}�
�C`H�th���5x��0ݥ��)B��U��d#��!gAI�RN�ԃhx-{n!�k�mE�I���Ͻ;��>i�>��ʸ����}p�g����������1M��3�gcB�<��۝�F7`_��h�DRʃ���Z���5�P���D�wY�@��U_��ȑ⮈�o�XlxVHYEB    fa00    1140���gF�������:CW�0�����oZ��'6Vg� W]�QU>�r}ZG%�c����G�u����,W����S�,Y��ʮ�����|}� ̼�?6�B���]�ѣ ��+�d� -�Nb����m�x
ɀ�~�7ې���g��X�&�eE0uh���/�S�^h?-EZ���a�jm��@Z^�X�@�.ω�h��i*O:j�p�k�A�,�1�40���z\�o����<��x����5�w��4�߂|��+ 	�6�������.���4��~)��G����|-hZ�K�����+巯�U6�����VO7h��x+oNYc;�9Y0����5�z�4�GV�\tD�z�2q}�6s���2��U�F��:^�{(^u�'����L���ɹ���	~gfm��6��t1�U���z����c�陡��{����� �]'�8�˥M�6�?���RQ0Y���x'|ݚ���|!�thL��7��~AE�%J�f�I��$���y�U�;~�3�@]�(/��{)�A���45�k�q.�ڳ`Ziά�f���{�;��m$#W�z4�[�
v��z:u�t
�����b1��y�Pj�,�#���K������96�8p��^�u*��º�(��j�N+f��R�v��*N��j�G���)�T#�}�9�l-c)QK�X��Odr��\��������1�Hl��`��\)���m�X��gΣ�9�L`��};Dǳ��)�wEZ�Ău���<[f�}���FN�*�qf��+пlN�EC���>��Glݘx�#��M������*B���#��@Q9牠�N~8κ��#\g��;_Z:��e�ڢ^��8�{���>�y���+�P��K�Z�aW6�����K����J�8^�-/2px� ���\�{� <)���lNkL)i��: �����&]��DOݝ�R��>ԝm8���7�+�}���~w�QԠb'��M�غ(��ۥ�愛Vv��#+ϱ��u���Յ��Πn��[.�|���f���J2!0&�sؖ�0h�>���`n��ܷ*�gf0f�e���8#��N�G���W�3��0��;����idӾZ�>�hc��ޝe������s�b>������g����G���I�v��x�㞊G؈�a�׿��aʯ������,,lX���E�su�#�v���}��N���	�@L�*V�y����Z�1'�FG�On�|X@��l�l�4�\��o���懷�p��,���g�v�A0DG��7yB�[MO�O��I5�0y}�s5�GRN�p,�*��t�$��$uL~�H�$ǝ^��9R�Xpџ�^�J�"�p����sW[K�o;�u����-m[<ٱ!^d����d)J��^����!p:p��z":|a�2�{/6t\�LF�ǀV��O���E�N�?OV�F{'�ܵ��o�(���j5���<Q�SK�Qv*P�7 �#�Ж� ���,s��O�<�홑%o}�UH��j����'f�@���v�WYL�ɶ���|ur#N����v%��C�vvX*5B���̥�9�'1��GB��Diە��V�X.� ��;�SR�д��T�
n�s,S%�����4��cFy]�cyG���1�c�?��Q���/U_w_7a�y��K�r zp�{���HuӴ~~<:G���J��]�����k�Ԟ.c/}�3� c�����[���L�y��#gO�"����:z��F���F��9v�g,4�yt���K����?�6w��C��G�lw.|`T˥�܊u|�H��|���/_��!vZ��Q��Zи��a��.���.jG-�@�����uH�΂�i1i�R,m#
��S(J�}|����B����o��!�ߞ�ʶW���\d �Tk�,�����+M���t񅾐0��|LBr���b�@�"|�um�ރ�sv�_4�JP1����s��������/�1�Ѷ��UP6��>t�G�_�5
�N�w�uf+���!U��w�wF�XQ��.�6��y�,ƳZ��5��>uvB��Eܰ�������{a� =��y�Q�fcA�uR�N�!�ѺJ})s&�o�R_��ׇT���L�KVw����s�vB�T�+�E\=RK��v�JF�V�ZN%����U$E����{OPH^���8�z�'��/�8�&�g�J o	��'x�m��,C��;K/�i�.��~�L��U�oί(��f[L8`����}��˻�nѱ=h͚�*s�*5��l��j��@鸎8�b��GXQ��c�|8��]72o��=�'pGH�(�^��z`�h@yK�n��J�3�F��I#W�n��AT��/���P�g4VW~����oו��ǰ�G-=��*Yfb��M�fW�6��3��|��!G��M=�dE�Ø'�-�3h�E�5`E�����KP�̵�g��2+�Z��Ej5A��g����rX&��gR\��%���)��Y��T�U�&Û��w�j������T�.S�s�<����h��dr���LG�6R]����ۜU��⼩m�t����;s���@�{<2��_P����K& �$/���3���7�-��<i±C0F�.v��xr����k��-���{�-0��?��w�ZFX����f�����B@^���Ԁ��~�ԹG!ͣ����h��'s��uq.�:�R�<��ǿHx�gF�c�$3�p�M���*���h<FFg"��R4�r~�����O���,�(w���,X(�g���6�&���d�mN"�e##V�̩�2!dp� u��͠qd�  g�G��1�����åi�R���ī�V�7�-�0);��U�93� ��ֽ�c�9t���]�Rǆ8�>A1�4�������KAti�%C��HD�p����<��f�;NXCgP~�%�:m�8��"t��N�凗R\պ�d��\��s3TH�A�;{�$M��|�>7�=�]�j�MqʞWp��6/&��E~���}����(˜���C�nRsP�=�L�1�6u��n�#��.����*J�t)n���fW�Y?f%ڿ���潛7)"�8��;IŔ���Bv���������n�����M�E��x�0_�E(��k]�ҤwLBa����sk4���f�J���F�@�~���l�vG�ƞ_Kd@T��3,�#���)皮��ܔL0�f�"<�"�_�7N7��f�|o 
�9��`q�r����+���MB[i�� �	�cQ�<����5�4�ח�E�e��"]�eg.�>�C de��^�q\F��N��KBP{��vuj��`�Mqp�5�MvF,�fqƶ�,�t}�L(#)WX�(f5O/�q���|mʌ�x��0��eA073�:�xb��)�Y��/��7J��Z��J���$`1!0qJ�	�ވg��G��\���}u-m9h|nƤ)�u���v���7W�[i[q[�L��9�8�؇���^^���OCE ^�mI+�F��CX�"U����<�z2�K��a�4ܽ_ƫ
8FeMQY��9�2\r緃�V�N���X�F�~��*a��/�����N��~��	'摻�B��-�32W�O��]�5L��MI��x�-%`�93�����秴��ۓ�S�/\\�:j�Q��(�z�x՞��D��,�zXĜgj+�ʝ�[�c���$��}����Hن�,�[HJXf2�4: ��p-%�?Cږ>H6�e;�v�=�����b����ŵ�c<I�\
_r2�[�֚�g�A*���G�zK��3Q)�D�T.� *�]ҥ���N�x���ߒv�5z�@��\I�?�	�O$zT1���=���{hCm�+��*�i��&\���v�sI�m���*ye��C�Y-b���Z�~h�h2ʣƄ\�N�0$�{3��#�������MW~��^Sq�|<��T�1A������*��=�V�=�݆RWl��)X�*Dћ�r���D�(�-�xg?2.&R�p5kC��x#����Bg�O��%F�J�0 J��[���2אJg (Gd����L��d.7U�`�H�����Aа��>��l�GV6pߗ/hr�ґQ�.h/ҌǍ%s�kIk�4�0�.VaMU��ZTg��e6Fw�X0����R.1��tG���R������a�C��{T�=���\`��}:�{T��Y a�a�N+ra�a��Xp�b6����p1-��N4뇸���':�i�w��f3���u��D9�$Ft�`P,�"BHp�y,����>jM�9~��PT��V��܃�l�{���
����f�mw?�}���I��v�gɷm��)�9�B��w�B�)�]� �6XlxVHYEB    fa00    12e0��8aF.�q��N����S4Xsb1h#��K�J�� :<�xzt~��z�������V���n��0��<��dT`�b�W�,��|O�0��q��(��I&s��z�:?v��BB��v��L����h���i>_�r<��!H���AE��ORnz�����lZC�� ��rZ�sN��-� ~;B ����k�W-a���*s(HEw=L���ף��a��[��ec��%�����@@��#�q�͂�LoLO��$0d{W��0b0���W�3�%�����x���-��f:���(C���d��W?��P�� �뛲��&o�
eJ�A���w�@��S!���3�o�Y�Ϙ#n��a7�g(��W �C6ݹ�K�U����a���aK90���hE�*d�����Nw6ɇ�{�F�9B5Z�UF�C�ǋ��4E�y��Yzo+���q���'L�(]�	�9���WG�����7��T.]gl��+��쀹Z����3\i�rsT�첻�J���4�6��Ub����ͫ�����iʈ]y�o��;6�J�~��J0��-L�l���#]qg�����u9���xkPX!g��gs��b&�p9�33gd�/���kO�a�zA&7�ox���HW2AaP�)��~��JI�97��6[8�]-�z��;���~�s��0k&��_�W�ѐ���UIS�aS�����2����#b%pR��y�쐸W���ÈJo��L�B���{��F�ŬdH��	�h���u;��a
���O�h:�;�1�������$��Vőqj�{)��-��!�Ұ�x�q�Q��X�"�#�@�0h����1�R��z]�(#�Ni����o�k4V�����竧���g��G�^�o�0,���� �v�٫NkQ��'�s�w���k�H��~
|++�T�-;�H>�u��8��W���m�Bp����	�&)v�6�f�;��	?���3���9Z?!�#�|(��,�]~��N*�p]���H9��|Q�h���'�!�4��,uT�Q*�=;����p�/�̲�hl��U����j �-a��!����L�#��a���|�%�-fW��zO������{�fڮ�N����`�sn��i�$�����-&�j�Q�2��am(�`��FR��r�v�����	O�}]S��WCsY���^�W�����I����N���hD���|���#v�B*��#��
`){�hwa���P�ӍFxI�����<���.�z�Ӭ����2}�H�A�A�M�k��D�B��Q�eL�����{�<���|�JV��xA��ab��]���O42OEi�g(h �Ăq�ɔxiL|Oc*�/��<é�X|M0��_ZP�P�j	E5!B�(W�CY��0�d������M�|���k�N��N؛9�~x,���u��	��� f_I6'�!�Qƃy0h$�}&��ap��<Q+�������lW�m>�Y
�0���l�%D%P�a,Cߔ �$������Ê�z��FyVZ	iH}��o^����FH߈!�&��z��6���Ü���d�y��K9{���;I�Q��2W�>� �1PcmGz�^���	� �qбN����S���)��h;�/j
�\��ߺM�;BqN���>g�(x�P+�M�j}E��4��K��e63
�b��&5B���
 ��5��V�Q��)����-�X�ET,�!{�:�(��U7���8�-7���,�Ӿ��N$P[N�F��QA��d�Pj�1��B7����P�e���c���&�B�2e}`�\�e_���Pd$i|������X���f)�V�~�>^�nRYrI�!P�ы*��N��{Q��o̋��ܮ6��6�5���<����2k�����t�dK-��Kk\藵;�@�7�}i�~� .v�I��-�G%8#F8�R1/���sy�ɩp!ZF��mI���oY߬9M�G:�I�op�ĳ}C,*j,q�}�X����V��Z���$e�"� 򘈞,�-�1�|�-ge��~���x��	K9Q{��s}�>;�ˢ�N��eᅧ�FGaR���W�5%��W�X����6W�8��v�z!5�k�?V��Eǋ����=�:E�O��`Ҹ�l=����I\ <l�xa�'�������7��l0�J)�8*�e��?&<Mmjd���M���F�rJ���*#v����GOS�r=5N&V��`���CF)�}Y��r}�jv.��)��am�ZS�QU���J5��\q�|4�+\#�/��&�4O�]�KV.0��(e]LL�il0��Gq��楪�=���)9�s���������:07R�c��=�C�4�U7��pB��oe�g֚��]�1,5����C�I��$ǉ��Mkk�6�C���ǘ���e�?40��y�5��?�c����0���+��ʘ���4U~%��.�9����]WE��˹&.M�c���=&r�9v��9U�U�|(��.�p���L�Ҽ`�
(�6�F�4���?�P9P��ДZf҃Ԕ���8���"_��AN^9aL����C<j��Htu�y�y��R;S>t׍�x`��P^��9�xV���/2XSt�ڬD�[��O@�%tɘv�&����Ƞ����'��|�	��x9*�����cm��k�'��q@A�;6�|q2l�'���@���Ⱒ$�:;�0X���=�͵�����:Y#κ���t}�Ъ���t�?#֤.���]�� G�4pMf[��yg�L�=�~dW�blXe	_ŭW90��B&�{��"��d�~�Π��*�!���Y%�е�@y��:lq�� �p�����KS�{�ێ���x)��hVK��y�RV��w��S���F
��ˠ
3g�r=`����±�����k�B�u;���-����RԜ'�^��C?n��_�3h8�/#}/EG��`���j�]����4���-1�yn0����_/�x�m&����k�Z��u4�[P�gۿ���G���2�����CޫF�ָ;���d]�X�?lϕ���8i��*���/�1�?�#kn�.�&�� -���9%�.e�W�ө���e���Ik�)�#�B��NS�#������I�KK�f�oˍJ��[6��٦��Gh8-'�jl�
�^���]��:�1��G�[h���?-'>�1П�̼%�U*\q�m���Y�{)����q�cL��q����\��XMB}�Ӌ�dҹ=�i�a�Q֧�W���ؕ:ʏ(�+5i
+ ��]`�A��Lc�����5�~�嶠���2V�[L�ZqL��W�`���Q�Y�Y���=���?{�O�깢�Rx;���N��S	�����=ˍ����7A2Z�7��>$A5��.���oS����*3�(ȦQvF���W��$���M2gh��Ƿ�t�5�($z&+h!�?#��\=��@�)�����Ͽ��j�)2rm��I�� �ޕ��m��?]'�<G�� iyQ�s쫈���2��/�;�=F��hzFN�d�W�+���.�K'6��Yo�H��ߴ���d�ޖ9��pL�t��!	u�ϩ
9.���hΝ��W�$t��$)s內��3$�Ҿ�l^:qglR#_��W1~���/��O\[�Lh����	��E<�8&�k����¢`2�d|8l0Т��\�G>߫��n�.6�����!Bj�p7��0X� �Śׄ�����3`h -�/��s�����3�P�V��ˏVN~Y���F����wW�u�vKvS�J�����l�I�,`��a��Z6G�WP��ʳ�Fƾ*K�G��i�K{��A��+đI�E���	���(���S�p��b<�7H0�@v� '��-��d�<8�ƣn�^
���0���_f�}&4�$�0CՁ$p��<���ٴ%�%=��&�"(\�Z�1�v\x"�R��@V}�z�w�ZNB/g�d��Z�$@�$'�K�N&��{Ԍe�q����m�P�;6���o�R���u�;RB�n�/�&���Zf���(V�	.�4�EC��KV;���)��7�9+�ڐ�B�`Y�J �b܏�k��g��M�X (��y:0>:��|��O��g��8���=1v�S����y�`Tr:��H�Dʁ�rB��p���Q$�� ��5��E*��& c�I��o�j�
��s!����"!*r)XO|*���Ϗo�Ŭ.����O�Lh3%���j�כGZSi7ӵ�N�)�#�G�$>0e(�c�ܾ�I�Rς�����E�@�r��� }^�YRh�7qF����w4K�*s�j}� �pZ�ќ��(xQ����>��7H�*��	`m�X�mb�T~��0�w	��Q�!+���P?&rWR�8�I�ə�� ;���3�3ޯ�Z&���/y�ԏe��u��_wFXsZ�?��솲:�I����h��J��>%]�Z�m��~G�<���%��$6A�o��{�T"�JeyK�@o���'K�/����MT}��M��Rg7��Ax[��)�#a�|)�Y�lcӸ`����EL)�Ms�iV��a �ܕ޿�g��!%Ag���
��ޏP����L+�X���T+��S3�[SLT�s����񕨏CS٘g�N9:�aJP���\k�K�!ɒy�ĉSSZ).+(?�,6�l��y��4*��2����Oގ���M13����2�4�ʽA��Dل�X�N���/�Wz��r�"����fl�2XlxVHYEB    fa00     f50E��v�R�z������rJ�s�������;���c��xp�)CϏ�g��$���b؀�	�Ag��s*�ۀ��GLb���)FPI�r#o>F��D����a�� �L��g�����-�L��EY���زN�՟�FE!�C� �y���?��s?�*�y����g����ْ<]� ��f����0�e�s R<ث=4#�dPX�&�Ԫr92ߟF�v��Wx�P��a�5����n�����n|�8�v��-QT���9|[v��f����������z�O��+cTn�Q��{e��F�K'�zߕt;�)8ǭ��a���Q3��R�������1�&���g��/��F�"�<�N��0#0/|��9H��g=꥖ї��Xo�o�:�&W">���B��N�!���E�����ݲudw4 �^��E�-��ոS�1�����W~�x=����Խ��Ƞ_8و�]���m�������diO Հ�H��tqq�ʒ�H�r|�ҡ�P ݪ�ӛf�|�,��+
��e�pH��=�X=��d�N>tE�}�6Z�'�/-�c\�F���8��p�MW���Fp�#v�ٮ��p�[�E��K���ul� :��ʲ9�X�Ql�+ n����懶��t�L����t6A��
�W`�3��8�b��cȥU�����䇬QAX
z���E�ج�Ƅo|�q�R�w��ܭқ?�o� �6Ƹ�p+�|������T��X2$����������� {44m��r�K�0��~~�������Z���:��7�O�ˡB�~83uf��LiBJ��� �綫J3]mq}������8��L���a��"G�d�L�fQ�����y���;2?�8�6h��]t#��6��'�����Č��TF�p��]��{oSJ��p���)L����U�	 �q:Е�',�l/�_V��@���ѠP�O��xf�\6��������Q,$����лP4�Pg����j����pҟG��W����#�ZOA����˿+^?��HB�#����(h��ν�n!��˒���9w��E^�ۊ�h��u��Z���U�H��y����#�Z�7aւKL���T�d!`��q��۵s��q�����k.U}�2���%���L#ֽ��}a�al�Ѝ�[Y �CC�H��=��~�M���:�:�^?Ր���AؾO�
��K�}Z�g��3��;�F���y���*���E���y��=(�l@�ܪ��/~�t��Ǟ+��Onľ5E��U�ٱ;�f�b�ɲ����H^{^͟�蘖Q<s*�Zg)2��ePNyGFQ+zdJ��<H �5�q3�K��wJ��7��@�Sz��.y����z-�D���]���(���.+�X`?��=a�a��.���gؐ7�?j��ɱcH'~��)�7S�%�hfO�&�i��Fn�)�1o1���D�R1��e�X Z��@�Z�4s3�ɤE\53@�;��iz����=�j��H���]��Sq�����i�[�"��ON�/6�	�;ZԸS̜*�l��Rl�թ�܂��Wy햎��绕9ɫ+z�6[�t����5[v�^e�"�"5:1�Q��&NW�_U�V���̏"ܳ׷"��\�+R|�\��"ȁ�X|�2A[����O:~���ǎ�A٨�+x�:5���\�F�璓�*q�tu�v�e�Y�������D ��g|� P�������)�g0�b�Ɣ�?P��I�����ɭ����8~�R����Z����h���A�b����?$���8'�kȱ�D�u�T�jt�Jo��2 �D������~�e�'*"�ᚮ z�62>����tVC�vh�Z�N��G�x6�$�����s�*K6R�KEOs��ʐ�Qc����a�͛Q��?��G�-݈�:l�A���������o�>��) M $"m�noc0�J���J����x24�y����5,�<��Ӟ V[��(������8���t)�p/8L���H�j�lٮ�n4���l�� �j�ԍ;®(��豍p��,�Wm~t�8E�6$1�=��G���2����󮦓w��
ƛ-j��r���l�ئIf㴉wSaR�,�^�Lq�����zL�zQ0��*����|����nҭ��_h�
�,��76��������_19�V�,lL��߬1�C��\�A�"2N����;�	�q�Mhf���=��=(��zӧW��x�7XكgNS!�uŎ����MC��-�E7�j��#�L��"�C�c݀��Ϯ�+�y��X�%�(e��GUC]m��/�lJ49L�_��~����%���yq�L��G��m�N?4�^��c�H<���:��Eo5�7��
�t#a��a?���Zף-�P�%�B�g6)n�5zM�^�q�}�+q
���k0��0�}7>N��̅&S`�M��?`��_�&;����T/��D�q��ve&���jYӁ��7D��RpbŎv�$�b-����v���qv|�k~ K"��]�/`أ+N|p��w���N�b��s�h��u��/=�
Z�#�3{����Z��a�V����y���ڜ67A�>e@��R" I߄ҵ��~idC�V�ی[Ք�<�j�
��H�CV��VH4ң�k���Yk�oK��H��ouv��y�k���
o��	q���.̐?��3��w"7{�n�b�VZH�y5@���W,ѧ�������?�P���jV��S��%4a\�ﮊ^Gn�J�w��߷�Z�~(��#.�7�/���
�(�L��K7���[�R;Q̤�,����?eSxb �%�.���փ a�A��`'�c�h���(�4�Gri��1d����Zqww�+�WC��gLp|���e�JN	�e��o�Ƒtf,�N���%e���fm>�{�Ok��h�K(ta+�����W�-�WB�r���踯�J��!f< �&����%�R:�o�I�\H�)�&���b/X&Z�/i�j�����F�̱O�k��/� +�� ��S�G.����C,��:���4>q?��Ϗښ&V��y�b�cf[+����A�W�����S ֺ�M�)^�c̕�wQJ���HA����pO��w�n?}��yp�k�LΣrl��~�R��!7@�

�`�޴�DJ�;$��f��σM,�����$��P�ް�M�4���N�2�2-�h�ᱷ���9�H��]&hw)���*������]~W:�����e�z^B�J��(��}{��p��FQ�>�Eiע�w�Av}~>�0������Q��-�xJ�����w��\腰�<�b�N<H�-;��i�����c	�t�U�r�݊�4y���j���ut�m���w�&gR-�%|O��z��)���X_i�@B���Q+�4A���É� ų��r�����Vw$z/#��?-F]���Dmi�x�lޟm##�7��u�8���:��g��:8A�u�6S��OeӒC&�����Ԇ��[KS�\.�N�κK�WW-��
�u��[��!�w�4�\d~N�ߜ	)�����;����!�~��������rި`i:����`�bS�.��1.��l�+g0E�d$��
�/U�`����|����E�w��#���ȄXd{���LW��h�6E�.�������|��ţ"3;�#�Jhk���mnW�V�\$G��!��%��*Rg�;r�KΞ�����t�b#J��~� /a̯�H���-�D}I�+yg�r����u��`�A��g�S���T���D5h�	Us�m���^~���FcH�>�R��Ѧ;咠s��Y*[�/����I�]�dY'r�-�<���z�)�:XlxVHYEB    7273     560h;n���2`���7��Q�w`2�%�D�&�9�*���ve!���D�ɇ��}���?��n���ӗ�lqN� �J=��u��<��f�<J�d5m+��u!�� 6Y��u���b�J��?��,��ś����Qq�v���5�v��p�M:G���S�u`��ɤ1��x���lĺ��a���ԅ�dRVq+�Q�[� [��|rr�L��%0�|�*��+-��G��p&�Yڈ)��|� �Vv}2%��f�%?�(O$glH-[���O��Oe���R6̖��Lf�� ����'e�����W _3;��Uzݩ����?�c��a�;�h~vâ�FÈV�<�ܼ)��ܖ�#��$�&L������͜��OGR6\�,���."�RoJ����Ԇ넒�qT<Tr��a�o!ʢ��qx{�[fA]�cz��ͭ��Z�d�K�9������H~j�YS��2K����;�����<�S\���u��4j����۴q6��7~�:�jY��S����B�m���(��	/�i�$▨.�����pX�:��eG؂��u�K�R�ߚ���:q\3�*L�]3��	�r�41�[�:���y�(��!2����og��.�{
Ԫ/�{�0z�)���ձ1vX���5DSP>�� 7/�*HDt.`)�~< z�D
RE�莋l�����]�B�2>��-��'dH1nG�m�0i<�����i01���&��7��A��cu�x�R_B�P�!�I���13Q�����I��v�v0Bm�F�] U��9y$��2��^�)����!��N���w�Lc�[�SP-��D�RJ�u�̎�p"
�2���[���
v���z�y����1���=ҭ�`�����5�AQ*o���
,���º��yV��O-��]��7:�#W�{����龂�!R�Gƛ|=cF�u�d����X`�!iɰL#me��	�.�6���� J� �@�te�!�ԍ5�џ���-״�|����R��:�������}V�R+��OK#�A%8/xPU��LM�_:�Or�Y#�� [z�.-0���:H���@N>�������w�d�C�a7݈��Dq�����VJ{�/�x��Ⱦ�q �aIq�n%Ž�֊ԦXI�C�"��)��3�����s���v6D@�|ܙ<�����S�DA�{)#�M��N��$��LՌ����O���RC�?��3����B�bǊ@-ͤ1���:樍��A�����e�:�f}�#���j0(�/���{�W΃84�*���s&�3T�w�2�g���H����K&ޝ��n�Ϩ���T��&�e^2� x�&�(�