XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����.�-��؉Wcu����s���V|�E�p�>i4ኦ�q����?I��7��e�'a��wQ��qC��-���*2hI��^�c�<������
�+�I��s�F�&�*_�	o�i�d�����=%�򋫪m,�E7��m�M��o�R����uoE����JOX-b�"S��~eѣr���-��^�^٘L�j���s/!Zp��H=_��+v#��b�C���\A�1�.E%8��Вj��nL>.��w�Qڟ�	�.�[ߪ���ა$�Fr�#�j���'��������h���z�����;��|��G�2�G�c��'��VS��y�(��YF��#b�_0F�Z�m�VEk��ٔـ��>XO���� g�-�����|�C�,��b���
���������<����ǋ��p�L���]S������r@��FR�e_.u�s�����7_�6*�m9)��]iug�2�Ʊ�ރ/�y�D���w��n$��R@ז�HB3��ytv
�
�HPYdFAp�Sx��l̤�zk��nt*���܅{�������Z�́�|2�^��ơ��Y�LH?,�j�1ͭa�8����4�����x��
anB��p����64�ør���1|�w�'� �����3��]j����2�_$m_�s����z�&�i ��@�R֗oEa��+W�jZ�`G�	 =��>4O�o���_���`1���F���k�����$�;LVn;^_R�"sm�XlxVHYEB    fa00    1fd0`E�L��y]:�Jp�l©Д���u�
'�8~�uU�}�5�rR���\z�$V�Oҟaxr�������O<�5@�|�8��[B�'[��&{RD,&\��LA࠿�����I؆��V�>�w��V����
9� � }%ٕ6�A�7o���@��}*D�/-]6�dJ����sK�=sl�L	��Au�b��:��Y\�c��Dk�--��i��}[oCNǘg�W��:�4�}���~��^�� f[E�xC ��}���cɮ��W�����\;�f�G�&|/��4s�G4D�.�O �:xC�c���E:"ؐnPL����"��o*�U�2�r�˲�!o�0�m~�W�ŎцC?��E�����>��\�x���D�ƻ�/�@%�F��˟:,���`0Η<ZqA�i1mp�g�}+Ks֠e�6�4ڷ3d*��C!O��%8`����j��o0��؝u�'ϊ��t��o0-���`� H���)�s!ՙ�¡%7��U�F ��c�������}��8!�b����ଁW�&W$��r���f
f������}W�3ZLUC������̊�p�x��a���٧�EE�����3��W5IY��|N�J5"3*�r�ï)�1U<&5c6�=a����W2Jlrb:����X]@r��GY�DTj(��bF��b#���V��1�}oea��x3�P4�CFr6��%������cx��a��S�XI9�(�J\��d-�P��]�� �^N�/3��@ى�&�̺2y�OwE���" �YCW^��Kp`Xqk��W���S$Kv~���}��4dۦ�"\#����Q�2�{j���M�hӒ�+)PI�;1����pSW�'KH�]�1����"k����=ȅ��D�[C�7����nB�P�R�9V��;����O���ƭ�'Q�ڌ��Pe�{�a����v�A����LǦ~��)m�'k���<�6��������:5�bS��T�c���>�.3�N�(A��O�0�Y�R��*ɋ]���R��M��g&V��"+�E�1d�o-����T��4U	a )v�R���� (Xϲg��8]7�ީ�[�js���=KB�]?ڙfwrt�YuB�d�h��&�7�a�m�h�)A����WY̫�۠vU���AB��{��]R�$OTɱ��L	$ο����d���B΃S�t�2sWߴ�$m&���#kP�,�10������^����fb�et�H�o������.�&l\3�K�H�*A��z~�w�x�ClU�6�s�ǻ�<{v��>J�\��O*v�i|b|q�˞��ΐ!U��^�ɠ�ؑ_�BK��I���4q�-�W�+�g�o�le�;��Jf�g2Qd�\�)G���芘�F�* k;���#���&S�Iݪ8�C��3vx`m4����qY:�{��c��K���|M��ʂ��5fq�;n.�����ܽf������<�~� |�M��n���5N^E�%�p�6;�.ݯ��I�C���f��L��\�l��M���㋴�1���5ƿ8Ҍg�^<�,˽�F�v���*$P��@ع��g9��%�V��v�wka����L�f .�2��򴺈�ARcR=�P��Dy�.W�I��G��lHm��Q6O'����,�wⷬR����Y(��-�����h7hҋ���ޥ��~�����K�����h�Pj!��J�6˺���J)��}8�J�n�!���,aDU8��֗��0\x�ᖺA��·ng�� ���P�q�ubJ*��e�۾���tA#���Sg=��a�=�|���aaP�	�R>�I�h�S��iT��F��?�AEm^��U��l1���=m�mS��J�na����81�c��\H��ՀP�V�,L9���G����J*T����;����6�w��r;��*�x��ƙ��9��T����$��]���Q��\Y`54��Qz�`����[/���U�A�\ӲZ�F�� �[�mn��.�4_�~
2�Tr���f����A���K�� �a��Aa�CV��U{%nu�p��7�ѥM�*�E����%DVb�U���f&ω�r������������I�7�ry��>��ܦ�L��M���GW�2�d�@�V�F���^�����#;A��,�)�e����ʷ�� $�}��*^z�_�]5| ?]�*l�=�Nǭ\`�D�?�;Ct�����«���j��Q���zr���6cHg��"�^b:L�#��ԧ�x��8hm��Cg^���>cr6Qm��;�T�0�;ES�f�.�|�p��!Q���pUP���T.-�k�ue��^ �?��E�X�SO��"�7�(]H���h1=m���&�J�9���#�9�{;F]�q�:s��l���ւ�I/���+�.��nX���f���	��������z$qg$�SW��0-美O��%�.N<�f-�;����7`�8�3�|�(���F��ܢ�$x��|"�.��KaR�~�b�L&{]��r<��\wQ����qB�����T;i8�?�o�B��!- �N�1�/����j%~]J�'�5?Ew��yO��N6^Qpz��7��5�Lk�q��A&}��g(�f1�1���H��n�@�A�A�zy���GQ�c7�����S��P�q�j"��dZ"��VJ�9d2�d�+�+��i�k�F[pv�*���էZ��L�	������2^F-��h��ӄb�*V����B���k�3nϙ�����}�3�\g_M������i��!3.����2��a�5.3��Ԣ��~�æ�wf��̹�ņl�쪡�A�f-�+�e7���Ә��x�)sǊh����޶ T&.{���}�t%��*��5��q����t�|
ʗ�s����C00)��ϔ�f������w`$�~�=/��,us�I#2��m�A����a��L���cnFu"AE}ZNR�^\�r�>����܁F�������s�)�v�?��DZ�ΧLvD����I�{X	72�d�5�`��B�	��B���H����b:�PQ�[�����o�UZ�C�*6���\�Մ��kg%�|��T&f#�p:IZ���X�9���z�y9���1�BubFSvFj��JDd�X9�!��#�zH���d!��Y�և�l��;�j�VbH�y-X,�2��1i���Cvb%�����PO��<Sg&��&s������0T��Z�j��6�Zl�
!$\�e��,�jR�0Ot�I����4vm�н�ى}=d�Ca�$�F��e�I��g�}L4Ej\�ߺ��ݽ��?����lbS9�E9���e�ҭc�����ׂc�꿬���q�0(Q��[3D��Պ���eW���_��qL~v.?�\�+���U������e �$YP������C|�(�)Q�7��E@)��u!�׉��i���!�q?jϖ�"�I�͓ACG&Ï��ȋ��hIF��j�8�y�z��J�Zj�Y[r������($�����	%�����:Z^|9�1`o#�#��u��7`�q��W��Z_�_:�	�ه����"iWƶ$2M�����r)e*�!�P�q��B����w�MP�5?�pE�w��'��R�z}������A�G��'�\0J3+{�M> ��G]����l0A�`O�
@��ň�{����cǭś�S �I�����9��
�SI�67��KU_��W�QC  �@1.�Zi��.�U�!q�,w��}Ja��c45yM��>8`��,t�����I���!�R��S!���'0	���uL��k����Z��|��8z����f�r��=��k�g�D� '��=�}��i�6� �B ���z����|�8a�8"����,��@J:�ې`�4�_~!����,�������g,E����;"�؃T��F��k�I`�z� �*�|̗�B���C�gT&e)�!�V�i�6����W�k�+~�c�d7s�߱a��T����2Q|�PXmA�$��R"���L��{����/�Hu�R��
�g=�V'���,�f�i����'O��}�929W��
������r=�<]�w�K}5@8�RK�� ���z�U��� ���9]|�ݒ t-�Qer�`&���tq����@���('�'b�=�u
;����S���M�KZr�yy��q?�N����uEm�N���$����X�= ��MB�51R�[Nu�F1d/%�����?�Q�"_b:GvX�z7B=�����7O�Z��X������ӥ�/"�I;�&/�͛�ŀ�X�^D�"�	v.\M��/��.~��Z��
�0������4��b��}�Q�)�4��vT��Ml:�b��!olJ0z�G{�Ό��hy�O����x��9�.��D:X���6�*�{������G`��a�9N-�Q[��_�=�=z�;s�OTi���.��'5�=���I[�L�����NJ�J�4H-.B.'�+��[�#�-H�x��S|�ծtI�/��/���skݫ"I�4#"���-� ? cǙ�.��dP���ub���d,��>Қh�K�(�_ـ��Ҋ�}�[�̬\ ��X�Cs�	�M`�rH�p#[�"��ɫE�<�}j�$�����f��A�����V����Y����[z|Z=2O��a������_�F���i�>b7��I���-~/hP��ܾ�&����oBf��F�vPr�g�2ijV�8c�G��� ��Io��ٖ��P)A��ٿ6m��fC�����Y���?Ʃ_`^j
b-���C�F.�G�U[z�扉��m�U:��A����XI��گ|\�C�ͦN*[�$F���R��D���/�����8@�RQ�����!u=h�q�$���Eҙ�[�`�q�H��.>��{(���$��,ʮ̾u��]rR�ϩ6�G�������4�W���K�e���L��Txު�~a)����CAY#gt�K���͓r-*�6�];yœ�1���&B��4ӥ��ur@�w�f1�o�x����ϹG�������X M�=�3rq��@��3C���V�|O'��ay�]����ٳ(���1�������o�J�2.���I�c�����(q;����$��hw�}��F_"R�bS
^:�RM���\,>>�0�ב����ؖL��r�\w��L�Ъ�T��>�C,-�7��%��,��U���9��b�?;aK���o��������jvs�]@�+���ó%ǮG�j/og����G�T!��. N�&Gb^dMI^���f�I�`����a&���-)7�~��ao�\Itt��d�8��6�2�n8�O*)�8�,��8�6T�R���|AeE!86��(�(�MƗA��נb'6C"_�ĖU~2��c��կQ�[nV�CTp�f~i�/��o�O:�d��.��}��.l�y�/8����I�?kW���]����3ܣ�1�E�0�}�@�{�dS(�ik��@Q�S����[W�z5�I�t�?~B�p)�m�e���H��-t�t8y�g8����#*0\��Y��Y�pB��X 0���&���L(U���?���@JғK���<j������
X
����Ji�W"��=]so���r|!���w.�}��3���o�����i*�/�9>'q�����QG�}fX����B>:�IE��w���	�?d���U�~�$p������>
��H��H}�����ѵ��qZ��W^��Ul�7/QH�a����l$�-��Z�����!1*�E��0�b��4i)�l�ގ3�>�	��.��F6Ar��]�#�ߋ	����G&��u���pG�>"3~�f�!�G
܇vc�!���-������)��U
�/��E��e��Ӑ�ql����hI�{�bW����b���H��9����������k͵,EhJ_ET����V?�J�0�G�PS9�n��W��ȋ��v�'�(J�{qΊ9x�c��j�:�[��)�~0X<*��nH�Z_�z�t�)҃Ev��Iu�?C9c�^P������!���8JH�7l'#Y�Ơ�w��/��Q`a��C�E��!��Ԕ�x��!I�hgdL���.�@+N$>�[O�G�\KEJ�;��Y�T9i�e�q�@�Zz��7|���"v ��_У5��욭pž�5r�8H�^9�H��.씦�֭p�-`��"G�H�iNN�?�63�6�=�,"�t�V��E���bY!r�q��b��x���&o"
Ka�<޽�-��*
.H򨆽b��΁J�,��5�l�����? ����'��c��|G��4�ë�C�!����g+H�je)���R��o�x � ���C:�Z�h/�ݥ&�vy@���941Y���?�#�N���T5�I�"1�'	U�6ƨ响phy�h��X�>���7��?%�܃<��JN�)5T��O1���2�ϤϜ�%تH����̦`����ĵ�M�����/�d�����L�\�!&��
��P����L��݇h�q����N�ͬM�3�� anj�����a�Ne���拸��PV�IcIHY�Qӱ��ơ�1��G�DK��'��򿚓�I�멼}.�R_䝚G��F���E�5Ĵ������^����*�	5#�R�پ�B��i�uy�I1�@۰r�����L�i���oV= �B�ni�<��A?��_5[�Is�>���a6�CKH{������E��7���� �:vZ�I�:zXA��#f�ǰ*�z���dG|�	2KU�����;J�歁�	��(/Hf�����=�V%�����Sϖbp�����jCy���%�f*P7�U(c�.�<�pMM�B:�y�E��b������If�L.g�heZ�޾{i0=�=n�����"�3&^9�H�0�Ǫ��Bפt��2軄� >�#J��%[��3�֒M���*���reN�j�D���4�} (~���,K��Zhwaf=��M��BL�?�������'�ցC�9��=����k�M�$��ZZ\��}l��^�u;�樘ꬿ��F��^�z`�W������C$�l��<��a���7㜼  �����gw����9l�Yh4\�Z���X�J3#�f��+'��s�=�r�t�'��S��|��M��@��1�j0�\�y�w�
��8/QJf3�}�~�M��'���}�D�@Y�&�ܞ��e<x�(��l	43z?ʉUh��ύh��,�u���*����(���ﱸ��<�F��$�*�
���B�k�2�;#i���G����UyWW���sX '�� �!cD���ѐ0ǽF�����m��9{���c����}r�c?Q�;�Ձ������gV��P|�1�j��6�t�bD�2�KE� �#�3B%{���-�!�9;����w.���+��J��K�ۀ �ѣ]�XF
܄�
�BZ��	�##z��}��gt�a:-ԍ���u�����#�n3�Q�_	n(��mω;����#��`BvlY�6��m٩Qd#��������|�_<�溄����To�Ӳ��������}��Ac4������9��V���'�Ma��kv?��	��G���Љ0y�H}��K#3OÜN����> �����ye����XԂ�bZ
�@;P�E��P��)�nX�Y��_�C��� or���;�k�5W{7 �,�/ �N�٨)�o���@)ۿ������Ik(�o6B�����<ǣ9�+낀�R��	s��^���v�UU2�+HO���h`�� u{��P�^Y�d����*��e#�{s`d���bR���ё�}�?�*�`c�L�ZS��"���d+ 0Vh���=�> q��U���<6bI��~��6���g^��Hk�Y��j�Z8�¹/�����qsZ%K��s�q���W�i`]�cf�I�	�bpQ�����^����jЯ�f�B8XlxVHYEB    fa00    1340�,\7!^���	l�V��Jf<DM�J��K�P�	�Z���<y�����;w��G+��J��p��n�5Ac��>_X�/F�c�i3>9��[�ܝ Yz�T⤘d��w��W2{�N��D�\3q ӂT2)KC�.Lu�69�:Y!��~�]�	�r��q�H_��Z�[a�6D�ś��,�ϧg�̓%�kj&V������?R����dá [�%Y����i�\k}ϱ$���� TlG"���9�8QZeZ�X<GCk,){e�i:>�v�}yx�2�&S�0o�|,Jf5�B���Ob���dg3/��#ɤ��{�)6$�*N�1���?Z���N�/n���n���s�jf�<���Jʴ�y-���ۂ�f����d3 ���2]�ݍL� E1[��M�iB�x�)�䗃��b�$;ߔ8�0e!6��='cg�4��a[� 7S��t���!8�魓�<%�C�k�c��[I�M�4ށƔ� ��F����$�X�Y��vo�1�k�Qx`\RO#�WҰR�DtWfS]��n��uB{�Yꉾ��Kx��i����Me���i��(���	lV��ʾ���<F�S1�����,�P��M�Ƴw���Pv9~I>�z�Ե;�f���X���vH��;p|;�h��."E+�5n��E&�;��|%g��.1<�ΡPT�5 +�l�u�!��>�DK:_�AI��jG{t.�A`"�k��fy>��
�o�����B�F�~�VS���"��h����M�-����wk���Q�@K­B��<���'������-3�w�g�|舋f��Hn���H��jhR%�ar��V���hK��ލ�	%\b�V���&�)�l�rĜ|���RJr,��h#��B�K�?�\?_W����?�24�?�p#tE�.Qܟ�2=�0Ϥ��% )�TuQ!B��8�,Q_5D\��t��M�ٿ���X|�/S麁 ��)sm�}N�j�'?'�^�TE��֡w>�!�'!���L(z+�w3�S����͘�0I`��h^��$��������[x7��F�Py��GT�������͙�M�[��C�	��j�!2h������
>��Ȟ�^ͳ�y�M,?�ϑ��B�pw[�Rccyp�1Q<h�wD[�Z�I�K9�o��q�dx'}�Vrp��&
�T՝��T��+X��N��F������D��v_ų���əDEmcڟ��ʐ�?��p��aº��G82�@��FS{����Ru��)8�Z��+��Z!��L"�<�AV�ݙ�O�1�+��28r7˾%�H!A��ف	:����=l��RӖ�3D�V�#��$,yS#V>T�~�p�G.�xFF��wʮ������Q�@�d�[js�&]���w^z�;�F�j��(�����{P��w$X>��=d������Ru<z�\�&}Θl��$�P���Z��'��HEc,3~���deDc��/��!�G�cRU����}����@1&�7}X�G�*�����8q*�����wp��#�~�D��!�ץC��Q�S��v��.I/`��ɬWzg�J�����
`�􏫕���w*��U�tO&�6vw� K}C�a���톚F�Y<F������|�QCpL��ʟ���S����Uf&S?h�ZU�mC�o�\�݀��YgB���U����u�w�|x�	��g�'Q����N�۴�&R��ڡ�g"r�Ǭ���[����G�l�c���HiX`7�+j oW�����c=�i4��r���"�vԻ�+���Wp4��"8hV�7�9NV��)����Hӕ��X��%N���aSq�TI�r����-Hr�!='�/��s�VA�2o�0�Q����Zf�D=��qlš4f�\o�AT��e ����F��.�'��+�l�7\}���mh$��������%�[������i��Q����+V��x�4]��'N�'��ns����U�����ltSֈ��7��6�/O2��U��5��A;��ۘ)�Eך1h�kҕ0'g� ���gP,Ո���,��s}T�r�z�~@�oި��h}\��meV�A> ��Ķ^�\F�,9F%�0��q�5��qX���}F���&u|��^�*(h���5QG�m��Y$���X��ڳҾK*V�S��dQ����GZ.����|MV��H�JM�z�F�����o�7�_}�Z�9�B0&�;�P��g���4��3�<�X�4��ց������0�u�tu �vz�ihO�}�m=�|i��X���+�q���@�Q��hU �Ǣv�9�q(V�(�,j�^��(X�?��ӡ�#�ו0pf�l��ې��)8�>j�ٹT	������T㭾VY'F�y<BU&�>�����k�y�Xc.oF`�S0&�8K^D[�ּN��WϷd��g퓎��Lʯ�2Qg���E���C������*(���޾(��i���:�b�����Ӕ�GV4�Xv�(��V/XPӤgQ'ز�A�9u��q��Ry���Ƙ#Q�$���&�h�o;���4���[�{��z�IJ�.6�6�L�M�54 -�"5~�i�l���x�v�:
��0��k�.%��m����!� jc��b��c��Z©� �˚~�"b��,�6��t+�n\��R�����4�NF�r�
x��`��}#:c�-��S���-K�\�9 ..v��T�r�|�I�zo�y�g�p�-ѿb��8�����#�]�)U���93VG
�ݼ��D�gK���"�ŉ�"7��e%�
�����/���|�m0�$�_�u�/��B-�p��/c�ޓ�b.�N�d�+D��̃.�4iߵ'��#��]�(O3P��%���EX���*9�e�����:�X'��[B��{�N� �;�$[��r"ϕ΁
08��0Rp�TV%o���<ni7I�g�?��ZQ>D
a���6Z��eyq�Vܐ[�-�����CE0GdD"�n="R{	�r�?L�{:hH�5�K�?�J��t+��*���7+������.�܄�+a[��f��(k/:�?�w��~��3��;��pL�Iu�t�̓��7��U��Ղ�;�e��3.ݤ��e/3�+&璋��2�Z�B�AL&8d����R�!�HA��L+�l2o4���5�W,~vzՂW�GC��:�!��5��%Chb36:qy= �mY�T��GG:V#|7�~v��I��Ȩ#�'���Ig�T��(�4?�JҬ�m1sg��e|�7��[dmt�#Sf����+>�{�l�w8#����I gc@A�]��:�X�_��"�Ҷ� |}𱑥�3��G���Z-��k�=�Ϧ���`?r�@2��_�=�LO\�2��=�=I��Tf$TY�Ş���8{�n�3�5�q^�9u��;>e	���e���w䱝{� PN�����7�/yz���[^�;�
�D�k?�+!ľ���?K�=@#��v�X�����/��E���ܫ�<������~!_j�#x�p�}[��tE�@=��GC��t&�z�����u���N\!��R,ɛ�/�u�+���Y>���ѩXS�j�ϼ7dO��$D�ǩ~bi,m��x������}16��s��l �~x�C��>�uṡ�4��T����@�*T�A��Ҭz�f�צ	G�����S�Ɣܓ�[�vp�9v�uI�=9��f+��������RR$�I�MI߮2�K+��^��5p�,�I�W�5�� !��Z����&�w�Y�Y�����qx4 ���]�v�⛕&����l�U���ϲ����$���i�����;���>����:��b�H�@n��r>#!�b>�kL]ȳ�{j����ԎШf��A��ڋ0��u�;�u{�����KӮ�2��eK��s'}�A��IEA��1�$ !f<�]��Q3���v��b����Bә帒#̴�_Rv�q�`�G��}0/�GHB��O�`׎ְ���B���lHx�J�c��BW>"7h�?%j�g����n�_5��� �Ү���'�^��f~q��8�lkw�j���9�������\�o�t�\O�w�+��Z�,�eC�kIT1�X��V8w7���EH�qd�2���pư��*e�j�V"KX�<�[���ׇnw���9�
��ܱ�_:ꟴ5"rP�� G6��z�?U�s�����J��#��3z\�$(��-�֙w:k!�@.]3CE������ଋ��j%2X�1n��k�ʃ��](NK&���ٸS:#Ft!�kG��A|�A%�?0��Q�ZSz#��������I�.&�se�S=���+cBr��7��N�b]�����#H0���\�m��4���*f.&R����D--p�G�CX^BϽTŬ��'��eHt*�;�;o���iD��,Ǧ�Q�֤=��g�檰*�KxG��9�hH+1��^�H)c�!�mG-�'�d�Y�]F�Z��|=������!���Rw$;���=E�()a�CĦp��c4Y�����n�R���$�d<�I�_X��ea�N��ۏ��{� 9y�cB��)%��J�)��
�ߜ�7<w�7�?�����w����r&��9FoP�Ý�ԉ����@��o�3��A���4"Ax���G�^uC���bUZ�y���H6I�����qN�@U�ϥ������*j^��ʒ�z�	S6ߕ�O�V�@'�HI��Q�m�<D�OQ**�8����I2C��E��\t�j*=£!��┛T �Y�d%LX_�-}EA85U�^ѥ�$L^��^�2.vu*�&4���g��B$X���p����w*����MpXlxVHYEB      e7      a0� +�~c�S� :*�ť�0�ƞT��0�6U� V{��u�eS��sק��z���z�Ա��ˑc�^j�W.�A�ۘ��jT$�GW�3 '��1���N,�\7s�1��W8�Y��Sǧ�+�F����ŝ���-m�3���Ba��U$�f���
�n