XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��s����X�&.b�F���	�rl�;�\��(ȉ��S�=*��^y�8�e$�T�<~tX�/�����޵K�]�ak�f�w����;�>�&fyl%��}�&��o̗$�bE$4�V%rC����k'u�_�`�ޟ<��zQ�c�Av���6�~��/3���H�?�|M�������p�"1ƌ�A�R2>���
�X�p��y�Ё���g���&�rm)v�F��\e�ɇ_����� \#Vdnx�a|>�m�!W]�n��^�I�c+�xjn�p�S��8�`�(R��E�q�R5��)�ۅ&��U~��VTb1�%l׷J���m�Ugc~��vQ��� �tp��mچb�����=q��o��R%Ӌ���[����w��H'�0o�+<jm>tW�����ZonY;��Lf��S��}M�&�d����_����m#V�����>���aN��_�/���?,p�Yp�g&��������m��:٢ތmLC D�?�ҿ�7;JA��X#3{�z{�� ���"MO���>���W(m�@��� ��@���<%�;r���3�,s�JL�
9\���[�(Aӧ�%5݆�m�V�I:2�wjg�(�A�����-ٛ��%���=�ku r"��8-����Ӳ�����ةr5^N@�h��5�fbC8�\�yC���cV��C��@ʏ�WUgwz9�WŒ����ڡ���ȭ�� ��]�쀜6�PIR����h�4,z6ĂP�O��.�%=g,XlxVHYEB    fa00    2520fYpd��Ij�'SY/�D�<�3��r��oĲFt7��p��D$��w�k���:..�h��QyZ���O;�-t�"�e4���� �<�e��F��ȏ���IPHt1x����ˆUK�L��I(X�M�})z����P�乍'��K_1�-������Y�Ғ��ԟ�|h�㭾hUM�g���%��Hn�'7��� ��]wUP�vJ ��5t���h��ol�0*�k_�3�_hl_0����J�~$ȍ(�����*�4.���:|�G��y/���T����G�l�1^$�)l�1�{L��;�� C�ΎFr`d�r���0�_�Q�zY�7?Vs�)_n�Ivϖ���Y1��t��U�CR�A�'C�dW�����=�!�� �w��u�����x��F�Y�V�I{��z�	̭�9�`�5�h��3�H��`Yc854#^��=K����{�O���2:��M������JC�֪S���I��0�Om�^��=��0&ǽ�I{��K5iZ
�n��1��&�@Us�0W��6S�No��n��+	jX�/�����آ/�ՆIS�)��C����d�EL✍b2țq�ƨlK92l$t�7��Y��/fG���0�A�h��r�"򳶰��Q7��c<LPLr�O��L�9'��]�o��?P.5Pb��j:�Q&O$�*%aˮ���n��<sU@<?g�2���pQI�(iOp��]�|�����z����v勠�e�r޵Bi'S�i5NI�ץ����f� �`>�Q��C�S�ĵ����ƈ���5f��J�����A�c�?NA��O퉕��/@lg/ѿ;������_��߃<NO�S�!~C\�B�����I�ൿuۄl^d6C-�S��?�[�Qp�L�
\����SVD|�I�`�l�'�q��h�}���G�����x�:%�Z[��B&����o��C1���ɺ���U��pk���K�U8��� ��X����|40���ȧo��8'�R����Z�ײ�vT^�Y��E���R�	k�ռ���Cqƭ�͙�s�m��V�b�1"8��d��x�*@�f�a��V4QB���7>��'B��.�����煗�aO�`�6y��r�Q(t$���	m�����w���f���Jݐ>i|]�6�5鲪ż�o�cT����%"�E�s�j�H��d��d��/v2��%��1Y�y��S�c���)����_W3NP�8� �ﺣ*�jA��<��]z@�Ց7��>����ާRb�7�����X(��:�����s�8�"+"����[�G�Jaa^�q�L*�
KhO/�S���W���>=��������_�w<�Z�������h�^�kN��&Ր��~z���`\�9�)�b��C��v,1L�W�W${�l^']�@��4�	$��n©�U�KD��:�D\:S��T�P3Em���\M8f�&�3͚��}ƫ�fZQ5�p[��4m7���Pгk�M��=��xPd=��L�CWf	�Z�񰰆�+2�t�5~����2�O�e�du]��M������}�z2,����O`�L���:�7��J�n�x�&`x��q�ך!�̣�g����5;���A>OF���&���r�����%o����}�I�0A(x��֠�uLւ��Q��=��Ǿ�$ϨT���k�}�'�j%���;��Y�J��;�G��2l�U�|U�g��"�� ��a̼t;KS0D�ͤ�l] ;F7M�Pp���v�x������L��b%ާ�MyVK"R}���
J${�&�Z�.յM�&�x��-}8�S�^�JY!�Qn�x�Fߩb|�ed���7hӢ�y�aNr���_�c�o�bl37"�G��xj��ðr��`
�Шw>��7@ĐA�ApqX�"���<2�����F�!3�M�x�\R�zbe"&nRl��מ���(&��A �M���ūP��M��Ih���R� �~������U�c{;�]���C�:6����������+=SQ��ɼ���l}q��3D����5#^F�}.�2�^��q��<�����s�f�o@��~��<��Xt�ʿ<Mm��� ����R�N���`�o����͈^��X�:ld��N����ଢ����<�|����X48��Y�����d���"�F�j�ܼT7�&�����67Γ��/�Pp��y��7k�Ş!�5x�Hh��zqq��`䄸� H+3�G�
��D�V��эM*[�k�[����]&fXޅ�t�Β�5�� R |�Ջ=!�D�/����au��<�V�H_>iD��F`ه��*<�W��*s �`m�`fE�gg��K�a��R��f�>�Ѝ�BLx��S�$�_EG��'�d�U��̚M�� ���R�n��OMnu!�^� ��/E.x��?��̭����|�l4��,��小ʇ#8�*������jJ�9�}�hHn�W.@PRF���) ]�o5�W�x7��O�(K�d ��-ݜ�K��lժq�4�����7|^�"v�n~x�=�݁�J�d���V���f:i��ѩIW��������m�w� -�=��>0&�İv�z��ؗ�e�����0:G�I�X���zD2s��>�7�^˲�Z ް���n]=Y��]̚i�ݽ`%�����{�K!!�oMx�;�p/�i�ZU��������~*�u�����_�*VG�*D��pt�彌O�|�0�!�l�i�u��m����׭��G�$¿ᔿoB��`<���^@�T�,�蔺P �j#�eD\�c����4S�M�|2���R��.ʨG�8��%�ٓg�j�����疥��!�I����w9�c�����}�^�@��!�E*_
�<�f��s��LGef���a���т.�`|��i���� -�T*
>�ط��2hY���"t<=z���;6�T0���ηLј��f� Zɒ5�F.��E�#�^���5�@��@Z`7�N�/`��h�#�|e�x*��`��By�mn�v	ʥ��p��^�w����"�R
�m��-�/�0��Aa�`���e��f�rM���ܐ@��Z*��q\mN54�O'	4��Ϳg��n�ý�ل��4"+�
�y��u��������[W�ftp􅥣{-��l���c�������WD�ű߰��� �n�&9�Ɔ�v�d�d? {�i�[?~�rr���%��&sQ?�]��s�Ss%<���>&QQg��p��U����P����.�����$��:��;����x/D��8\+X�;CH<)ds�ؚ��6�T�[�� 剗
πA���$/�@Ũ��eL��۝<e�ƒ{DσY�O��x�a��O�<�m(-ӹY�������K�m�����c�*W��� 7��UG@�ZW��2���lh�w��Oر�@��|��zd��!6��2�$�����;��V!��{�nb]!� �0�8A�{�ԢB�vH�i��M�rlb�y������ll�&�$Y�P�.�@}�	���s�i��D�6��J�O�r6��r������@�Xd^�cB����p+�����m��5ӔEQ�+�<���ZQ��H<3�EH��,9�j	q�J~�d�f�f�~�1��0St��p�!.�{e�b�d�C�#ߚU��k
#]���~�#���y;��Ê�A���Ё>멆�{��1�685#~��������=R\ 8���p�1�BO�7Py���(�f0X���!#��5]��YdLUL��P��3�_��z0L�!W��)%C�ɬ�^��=�Zۈx�6�����>G͆�Ý��"\�H��\h�b�#{���{��5\�(ޠ�R�5 �`#�� ������/�.!�PF.�������j�R�y��sK�~+`ĩV�	[������O��Q�I�ڧ�z�� zB��b����w�\]M���f4\~z�ٌ.x5�c&k	u{Sw"�4IO�Y۸/��v^7ԺWs�T]E,d�Μ[�9;aI�-������ܖI~� �ѴX�$
��"a�S�Mq�7=�z�8��Af�}8\��|�Б����-l��{����F=�C��a�EDGdQ|�7���kp���.���4Ρ�j�o?�A>��0U�j�r�jx	��m�1*��jB������E,Q����}�S���i!+����pA.�&��_U��l4�Գo)[�mد���$#2��?!�YV�SP��>��O}8�P$=�7*��BS �a��@�
�?��B�縩le�gXc wr�i��(��W�a�ʶ��z�a�,��n,�E�� �8�v��P���/+�%v��Ts�Gqm�Uŵ����0��Y,�oI���@ӱ�
y\UT7F+�t�?���diz�C��62��oX��*0h�,b�ıs���X 8�3~0�&/�0�i�P���J��9�m,ͫ�gZ0�5pǎ
��zƟح�+ES,%G���):�?��ܘ����9.�%���Ol�� g
;#ɹl�!wɑ��}-nȨ*�*�����Q���0v�^�a���2#��  H3bԄ!��l�>[��8R�:~;�a�(�إ�]JK�+��J�P7Yq*F�!��垌a������/5�8ܠSuJ���UJGS�>�\Oc�S\i�穱��\����[�������!�O�Z�~�Z������Q���Ǡ����T�Meo� WVJlMvqS!_�F�4���~/�4ݿ�fmw��	J��� �Y��ħ{�w�כ߼rU�q��ȊO�cM��S���~}`:�>#D�]�JN��Z/�Ǝ�[��
Ӯ�ي ��uY���O�2�$3���\6��*����)������]�H�!�k�A�]�1�& m�h�j��?�X͒6Z� ���a�����>aQ��>�lz˗�Ł2 ��] v(p���,���w�m�G㯪�?v��"��k�0�m���i�c�tL�~�� O�VO�=���>�#�t���fk���*i���3D-��_Mya�W��1E�f�RЕ���]�;�hR6��؍��� ]�vU�/C꼅_����y[�w ��b�&.�6�7z[<.Q�ź|mpc�w��[��N\Z�v.G�����v|�U>������h��f'��;�%���!�{��;��6�1��1)Μ�X��$�ӟ�1��1���t�@��Ϝ2�l�b�����	���ګ�54�7V�߱���^�|T�e�l`dr�Q�;Ȕz|�WA�Z��^�I���-�e���8�����Аkj2�Z�~v��:�)>���z�z���J��oVĽ�c)T,��Q^ӿk $��C���ƛ��4��A?nS�KN�l������9M����Zߏ��K���d��g4i(H_V��\���PB�������+8{�2n%�d�~���?�p%R����h�V���%�(~����h��6���x �x�����69"��|�#����֢�
QN8_D��R3f���n��=5w��(!�8z�m��!(8�i2 ��{zKr�	�g�JV~[��}J����:� ��4��:8����>�+�_9V�iu"6[�ۙ!�0Uǁ���j�j�qm*�0K�|��c�_�i���&�zS&4��	�����Qv����]mZ��ǔ>?�{0�0Wm2yZW��'�wV������nԮ%�ݕ�'� aϲ1C��h��Q��#FOޣsR�e3�!s�?Y����$�l��ޞF���/k��-��M�$]��zƒ�+i�`�4�j�����ϕ}F@���$�c�ƅ��϶�F����W�´s6mS��Ʈ����������n�~ik��Cf��1���ǂV�����֝w80���x���F��I,��{�T05�������J���7�������[�,�� ��\X,��h5�F�d�����W-��I��]�`�1+���@�Kmo�.[n� �q�˧���~��`�qnS�$"� ���,�����m��	�����}�zM�.�r���#�4'���t�������ڱ�̢.1����(�X#���t�Oiwm�m��%�:�+�U��S<�n.��m�h�V���C",��(g��쨰��o �͇zql>P�فo�螞��HU C�om0K���e|{�����L��y���.�j�7���C���*���+��Ax�6�����`Y���N��
_l���7�,g��t3n��q��K���*���`SE�^nn_K[�v�y+ҏ�su-Bo[�����D:�ԁ����rk<Ck�%��K��OyO�xg�,���s�R��l�xվOK�ڡ���b �m�)�5[��.ưs��Cd�J���j� �P�}L�PI�L,����_���.�Ϡv���֍Ht�:�Hc
�`�6����8kk�(�Qp���=k��z��LC��o'�~�XɁie9XU%�=�[���wO+؛k� �,��-�R�j;�ܟ��g�P�Qfr3R.�ʯDY:�m�r7�ȅ�a,{����]A�'A`Q�,�V�^�A�cY��}zR�K+��Ÿ��m+�-8�Α�W䁁ƺG����|��/��/����NNH-�MHiN�L��$q�\�h�
�*֛0��s��
��p����Ӽ��b�0^iE�¬VE�6��[y�S1N�����Xи�7n�q"�\-(.��b���>.���-$N���LWm�_���[pi<R՝�C��TN�Nq[R'�:q�NAr� ���Jw�?`V�tb0x_��pX�EI(J2��*R��l�f�
1P �� f垯����8���mh����Ts����*0b�O��V �Ż^�P��ͮۅ�\O%��/�a<0�RE�IN�2EV,W-��T�VB}[��c��)�nש2��Xw&XX�Ppʛ������1��,��D7��Phti ���Z�+�aC�Ǔ��څ��9�RsR^� @�a��L��������0��]�¡�y�7��4���.�L�( ��K��*�|r�}^C�}V�����[����;�K@��%y��v�|fÓ`��u��,:���Q�L�� #R����>�.YS�>�2]�m�>fQ�P�J�U��*�EX4��xx�H�!8�!�y��7Tf�{��_�����<)KM$X�%�`��ory�"W˯l�u��}�>�|_�[`m����ceչ�F��m<Ѱò����q�`�BLGO�H
+�k��H&�d_�d�Ք/�3p>���qv86���[�fZ�;��Jo+>�E�J�JP1���� ɐ�kS7:�R�qE�
&�Cf�
7q����3"L���s����{^Q\/(ҏ�$�(�pm�@�x���%�I��ɇ�.���������E��̅�Ot����@���)|�I{�~�����A�s���%���m�|�����|#U ����	�l_�7���:���
�><��qQRV�ur,��$�O�D��kl�4Q���E�I�k���Dh�z�c���N��\ ac���7s��YhKP��EN�>�,�8�t�Z+�B�ܹ#�{Fr�l���ן�����~����ط��@+)�`�?dg���Z���=h�iq,0qݵd7��~>M��\�&�++ ����f�HrM�$0���|�/�Ӈ*����ڒ�w-����rx��l6t��� T��\��cйlV�~,������0����u��K���*��3�.�"[r����oR#��7gt�5"ט��֨��s��b�7Y6�S�,mwf�Tdf?�
b��1��b�&��E�!hw.������i@m��1e��U��l������qǲ.2�C���\�DގI}6�M)Gs)<��.p�+~��!��,��"4����9���b�����,.��72���Th�Ş��������{?�F=��&�3L���wp!'OY^`�_��	{��K�~�թ�c�k�6]ً�������I{~�%�O�q8�t M����!��!�W�u^f�Ib��r�WoҤ�ʶ9�5��=�ً y/�nIuWݐ�����]<?�C��-�T��w�|�W��7�(ۣ�6��7p��w,z�b�@���3����֐h��B��r2#�}Lw�"r��M)����d�5>�u����S���Y��-�R��l^�T�z��������~�qJXLr6m�����d���d���rr@Ӯ�v6M���ε-���%=Ķw���V�@p���ڽ��H��q�}�̶�qX�j�ߝ�_"!�(��r�1DegB����v�R��o��<oja��=���$���,�r*�P��8�ۻ�!��u��[(��sp�JƠYr������p�LB�ՂN�-���
 �4�:2g귞�&�?�!��
:��Ș��-ʻ���G������4P#]Q�k�j8�ϞM X85s��n^�%�(�L�	����sW�#�-��D�b�W#��_	�,Q��,�-���ݧ�y����0 3�|Hb���/&�q]]Nt�V7��x� ���C|i�-|��{Y�����g6�Ѭ��8������J���4�x��bA�D�x�����R����xΝsJ5U�~���i�ß(Ȗa	���\�2�7s�-�}»�5����aJm���(&�Bz�QT�{W>v�n��.U7	��;�z�]�u��:��US����R0� {dmSp}3&QC�Q����p��Pvx���FY68��/e�`5�Q�H@��(�Ǳ������L��*�����V��wh�"��{�����~*�ЈlˈT��(sD�JM�����X�s_u/bS#���z����$"�VbP�tfm�_37�-��JK<�%�K�yD�I�^7iT�uHz���� )����w��f�����к�y�+ѡ���=gP�Y٘�t7���+���Td�!"6�@���`1:[�����խ�P���L�����揷�A��T�1�ۅc;8�L��z�cBV�6\�0�w!�26���+�E6�P��>���.ExA�Ќ���K\����*Y@��� �&��ٍp$J�fΘ~�MH�|�Un�bH�df� �T���A�^�����v��f:pJ�Ȧ�A͵�N����i�@!��uM3�d��|�����}|�����h�?��}��������gɡ�6�bJ�e���i��4���߉���.�0���t�"��Jm��Y�4 a�6��<5Hk���²�3��V��cGz�=%-��|�w�.���S�\џ�3>è�(~���=��7�^HN�3(<�Em@!}��Sk�SC6�FA�o�z�kN��v"��[_� �!*��y�L�XlxVHYEB    fa00    13e0/��`��ͅG+�� |@�(��G�?X:�D����}�0�<�h)Q0��P{wEz18/8��7�����$����D"x�t2�ۛ�$&�D�V���tn[:��m'M��$���s��}��Gk�fc:���z˝��KD�,~W369�{�����zPɨ51ۥ���=��]��T�L��e!�/��C�لA��3&>`��p7�A6:���T~�����5z8�'ng[�ǆI�^d��4�r�7�"d��G��ڡ�$��`I{���xݺ��SaG��՘6�\TU������zň��ux-��Ћ��s`6̂�d�̥���T�à6���OC�cyz�~�<{q�[!f�"��0s~V��l�p�\�ޫ���[j�p�v��[�3俺�~+T���CC��
�1-0�y
6g��k��^F-�.���~���뷲��$*@�wӦ)����	](9����S�{J�z��'	�v��r6�K�t)@Ѩ#h��V�A�欼�}T��\���B�6��a���o�땀�S��1��`����ϲ��l��Ś��.~�v�޶4+�����,&���ʅ�TqfAf3U���E!���bT��?b� �p���|�oS��h�&X��(x�#~��B���>.0`��1ޔ�e�7Z��鴰�;�c��֣� jk3����s����K9�XM%7p�N���y����S���
&,s@�]���MB#���&�?����5Y��y1�[4�ML�`���FB�8I�L%A�mz�uߟ�PjݶL�0�s�\E>`|&�����jMͤH�����)B9)r+ ���V������P��=+���q�L���)������_��z\�m۹�ڃ��:C�s,�ԣ�?І�޺���Jc�вٷ�9��	i~��.q�>��P0��@Qer��@�ZB����1��9��ݘ%{��#8�Ss�g�%��T��K"kBEKA
�̵�K����l!4�h�/Zc|���4��4	z]y�b�2�8z�"׹Ԍo`R���n��shZ 3~�:�W�J�-��ڪ�~�!,#�);�D�a�1�`G@��6�XA����˥��V/W��� �͘|Z.�~��U����b�����{p�0�EVl�Bf,�P�,�Z�v�jοxf[�_���|�@�l�6F�Η5AprW���ͧ�O�^9ї��Ԑ<�u��"����B�բ�l��on27�]C��x��<Z[ K�B�@wB�u�q��q�8������)���L� �T�&�:�t�3�<�j �^��VS$N�Z�6_WB#�!��/-���+�r��C_k*h��i�f�/�{ϫ��I��dӺް%7��)�\^�Hf���R�TF�b��r�D����Y'��n- ۮEٳ�1?��+�vj�D?�]��u��Ð#��~o9I����vE��,9��}�wG3�i,>����.I^��]��� 0bF^eT`.���C�;%}��2Sˈ���%\����<!��x:A]b�#o�<��LoY�;a�qF�W���t�c�E�JnL��2y���̶vv�Dj-H��%��H����,�xOk��k-»bt�r����w��Y�'�%Z7@@_Ј��1�!?�`��G|��v&SS!K�žD.l"3@�B*{�6G)��`��Hb�OH]ԝg��k��1Ϟ��ɡDR�j(K�t��6��*�JA���<�+�#[}�A�t��\a��o;|��+@�����t�[��
����0�߲���HJ;נ��Z��͞�~T��xd,(�@>
Ti�	U�pBe�t�6���Lc�6=5w�����G��jJ�� �;�P�`�f|9� z��vl.�M7����zH±H��G��_��#,R���o����>�XP�8�֪t�&Z"��hSt9�a����u^�2��k�SO5����-�>$�������+��@MS���vvZmvY'�wk1�F�cʺ�YJ*����[��>[�^�u�D]�g�����i���ܳ��fG�%8/�o��{pS���ǆ@0�0"$u�$��4/K��$!'G7{xR���u� N\������ ��Z�wP�6��X>26����Uk��1.R5p�/y.l>�Q@�|�U�A1�LK��=�f`͋X���ŠH�F��%�-kU��so�1$-�f2��Q
����H5ː7�K�F��[�&4߄��5�R9�'s�~	�7MDL#��(2��h�:�5��pƎϰ��"�����5��h����F�iu�O>@���M=Z�Iz2H|��om�vO�%��&f�B ��6�M��ʊ�����<���m�f����6T����ă&]���p���:,���pd�D�ly��3j�yT� �R��8�rUL�E!�b��!!�����b{��5��o"=�BҜ�{ȸ�K.�g+:ߣ)��B:ܤ��}��"K�(UQr@F����yAu�����3�	h�K�91��M�5�,�"]��V8���7�����D5j�ږ�m`�g��۪#&�zsṯ�p]�Fa)�S����\�5�mt���-�$'��Pe��1��.E:w�[)��.�D7@X]�z��u���@�Ya!�P��,	��-G���زw�r��ǐj$��=D�P*��<m63���}��U��QL�R4r\��J5Q���N1	͝���n������E���?���cJ%ݭ�|�O��h�/�;$4��9pa�2U
z�p#{���%g�����ޱ���ݤд��i��톻�kx������v��d�h^o����9���ȉ� �� �Y�ؾZh�'TNfX/Qc��6�(�3�d�g�ȟ����.ѝ;���B�s�gFI�����aQW\�[j6��Y���8d{����i�/DKI�m�����՗����at���D����%�yf�f�7y#���\�J���qN�/�Õ��QJ��ҧT�����x�PP"���<8��j�z�����k�$���n��eD��~�ԅ���5�?���K&z�Z莏�����d���o���AC��������X�9�J�zhz[V9��2�NJAs�o�;�L�¹�����o��k�q��r��W!w	�&�����;����Fo��$�D��!�`���R�ʋ�iԣ��b�eދ��:��������' ;V*J��=��=h�Kf\�>�y]I�]S��R�*0�6�I��bF�I}	��k sit(�_B�F�=�������AK�;���	���ro��C�;b*����)q�K���-��/���{�����)�no ����bBxS2�Ѵj��|]j9h�n$� ��j�b �f�\����k�@��������PKu1���#�/N�[
("(��_0���<�`|�j�q�c�Ԑ�,����W8��,ޱ5�Ќ�k��.T�+��Q6��0NL�t�v&+D���^K��qy�c��{�)���"a��ڵ��ᅰi�4�r��o�zq��n�?��%��N�JX�nD������ӑWP�Rn}6D!ު�Љ��p��9ًȝ�ܵG.`G6��� ����nWm{a�<']��P�k�Fʰ��|�/��~$+گ)�u֎c�ɘq�������ku˥�M9ɉ�<ٻW6��h
1Qȸ�x���ϣ�Hr֟�@DS�'���e�{?$��b)��X�8D��&��� K%b�\��4�g$?�e���Yt�zw�j��#A�5�p磤�	�7���3!������U`/=��N�� L�=V��D��%R5���z�<k�j^�g㱏*җ��i��Q*�U���(��8U�._���4����\��Ek.b>G�bB���b�u �-���q �E�unHc�~���-�t�\���( 6�O��i:nF�V��}xy������"�4M�폵5H<;5�,��ɗ�,��og�u$&
K��u����5`�[߇�G�V�q����M����%[�<L��=�ۊ{��6�*1�b���*�I�	�p�L+C�A���(j��>k$���>)�9��=J,�|�u�w��zI�����@M���l#�_gb�/��b%��7����R�Yd�����C�'�8gD�g)jh�s��Ӹ��� �[��/
���� ��P��l�t�;�u�N�迉&�xd�馫����2-��/l�$C�����>�Q�*�=�vv~�'�\h8�u}�3wn���Js�; 1i0��Ei^��l坏sz������' P3r@,�����F�>#�)�\Q�J��KL篐�uu<�Yʞ�Y6jo����t���!a1�ԅa敻��#�*|\o^��A�w�x�4�5wM5�:�љj����B8�]I�U֡��Tk�P׽�zI�19�bR@}���T�{��@�M� 6S˽�h���q�j��ݙ�1y��8d��g��W������hW�ά9c^~��V�����ʎkt�϶4��x~���;�P�Rfu�+�3w��Zj�";U}���%�6HW-p��*X�1xG��XY�m��������Dkg��s�u�����ƥ�)��"5sq�n���r����_0�����
Eٺ���L�]l߹V?�8ҫ�S4⏴l���ͮs�E���Ѯ_�<g�D��S�"�v����L�+���H�e��z�ec!����Z�3a�(�9WTX��`j�9������a�iV��V�t�/�?A�o��S0���M�Z
jcb@'��>��["/���Km����[b}~�|�w
���s�5���W`-�MBݥ�`��L&�L$���P�2�K�ـˇ�Ul��y/���"<�,�fE	��pԇ?t�br+w�lD� � M�L(n��8
�ڳ�����'ShK\�l�#r�d�����r���¨7�vu{�bw� ,Nl�S��FB���b����Lw���H����bQɞ|�_�#�Յ���X�Z�uG�G���)���S� �g�C45pG�$t���Y�cUr���m�0R�x�h�R\�%Ĉ�AQ�TP⪙�jq�<ʇ9��w['�>b��XlxVHYEB    fa00    1780��۫�=�_���q��h(���D�����������pP�Hߞn�[�ӭ�D/ʆB�����S�����������wQ�n|�$n���aJ\I^1n)�EG�̚�I��D���@��xh@ڔ�2ȵH�?cr���ո�%��%c��ze'D�.9��\JEQw -�hLi��<���T��j��Be��� *Kz���"��]�ӐR/�p��uc1Br��f`^�S�K��h��:ӳ߻��0b�*x��ˋhN���WP�D�i��Q_]:#��	kf#Gښ�d��8�x����{(��2^q�����*�_���Ub̕���Gw�e����D�j�Xk�ܸ����q7�j]�� /���'|1*�#�,�35O~P�1i%���G�4�.Ҹ �h;¨Kg!(#VWm�v��ajx��ƃ,�Y�p�9��΢��E���'���2��ۻ���ׂY��F���Z�^f�@�����W��{�����6�5yjz<>#��yp��f�'��µXZ��w4b~��E��MM/��CE�ϖ��9 -�3�i͓��q����h�g�6"tA&�Ӥ��
��3L,�
~�32��9OQ|>�@�� �`>��:��Kgs_"��D?��+�Q+s0�A�	t�Y��ha&!>G����wڿ����6Lt����,����!�ѕ������*ϙ��aE\��h�):��cN!��5 �����V'��lf����ELg��ݧ�05Ɍ�]�!���1�3�,�?;!�^a%k[�W֓Wz�@���JxK���Hh�2���bM:�,�h��,-	�SN�K �nTf����xT2�a�Y�.��� ����&��πE_���B��!e[O�Ҕ�Ѐ3*�Y��=U�!d�y�g�4��:A�,.���e��(�Δ ݳ�b��~�Q�$�*6�����>و���"ï�z��U�/;
�Dvj�p��~�^#�Q�۫-��+7�엞�|NE]�?S�k/	�$/�j���YM'\,�� Z��H>�
���NY76 ��M}�'�]>,^��z�Bj'��B���	x ��4��q-�o�=�X�hh{Ɛ�I���ybC�� ��
Zi�6n��&��b������.l�3ϐh蘑\���;�޿[j���5}/���`6gV�$ۻ�AI�q�Z .���5m�a�)۩A���<&T�@5�"��K��ꮵ��͔��j��2�l�<�VT{�8J���A��I��,�+����|�9�y�i��&*�>j]�=O�ZJ��d#B|x��"��������M$p�G��/�};E�eά�&Xω�L�j�#\]�����v����)h6RC��7-��g��@ry��C�+�]�V-��8�"T��H,�^Ii7���HZ���r������q��� M��L	��>}�_{��U�~�Lq�{Y �Zr��caCKS�����z[��J���<��f��P}$������d�&��Q��c"�������禬X{wQS�dZ�FW��mX.��&P7�c�6]@�n���2Y����,q;�SW�v��/@B�N��߯�.*[VKmt� X�����c��R�,f�,����8�A��xmމ�,5%��B��%l�S�b�|�@�]w�C�l���?����q4^G��p�`�9�<���LZ$�]%��e�tM�\�147J�_��4M�`mk���r����CG.nv�V�6���~ˉe�tec��LF��\P^�Z��ja�VR{v��N�3Ϡ+c�@{9�I8-7�s�`rO)OE���1ܫ,:IX�_-��{�R�yS]%M���}�IQ8}|����}�@!7ꮁ���U�h7Ft�7nq4@-t�_����[��?`.�4�eN�{^��� |����J���$_�Y�4U@��93��/���ݕ�[�'��: �)����(�`3������-�h��I,�l�Nk�w]�	�8�L����zQЙ��F�P"J2�ȑ*��ʥ�q�hy禹�z!g�}�(�$���sT(>J���
2%�gy[�Т0�q8��GK���;��fY*i���Ng^�<�����19C��`A��G��6+�`���˹t�f�io[:�T�+���'U����%��n�3�$P��d���'u'Z��m�;xg�nt� Z�LsO��о�hϠ��8�� ׇRK�[������������1�q���@��R����^�C��[5@���a-��Ȼ#��]��uq����&���U"�ZX�Λ �����"A4��	��$9�^E}��:�fnwr�C$W95=(������ƅ�`�Uu:��˳B7��߾���pTc�Y�Y
(Ϩ��~�6�/��5$G#����N����)W x8����)g�j�S[�����lo���G��}�л��;�Y[�v뮵�~���6V�f�ޮ!�엌�'f���ǧ�.RQ�@�x�w_��(P3��UR^C�c��X���0�,���]��HE�/�)�s����D;A3
�^+�\r�f RU���b�s�H��Ys�$a&\��j��q�z�r������$��MU@�|[i1�9ko��2@�#wdc)T�`��8 >D4�ކ�m�C�U+�o�V��_�׆$_���uO����A�Y���
�7Pi��q{�<����t�ZQ�Ԕ�U�]����U4J�lZM*o�?f��J}���[l�3~t�DO�nɜ#K�>��T��y�;  ��[���-��Rբ�6����jI[j�/P�H}��d��d��+K��mX��%!n���/����q��1��,��R�vI_Gb��,h���q���V?/�R�/�sVÚK�;s+w`�� )p0������dĪ���������M���|q�[\\R�p)G��[�]$1ה_]��N9/�c�	3J�Lm&�{�lK��a$U��!,a9��n��Dh���jƅM��aP�����=���#hĦR��Brh��1�t:��
(��kL������²Pc\h�P)ըnj�G��ͥ����|�q��~5��򺆹Nߊ�g�v����Q_W6��ov�\�,�]�s�L~J�'[�ғ���h2($"����m���BH��uq�[���-_��TAE�r��=K����r66� ��;t[��uM���:�'z�w���'�kO���F}�wv�ֹp��c��=�yt������6�¿P���8�қ�78v�In�ܘ� �-`m�*���}_�F{C��"0l���\�����(e�c�oE ��g���=U�Ӧ.IԽ�V��I�Q�i����z0�ƃ�^��X�Nd4�* �E�tT]f5�����7^�IV6q8@�h��8]���\O�"�rk�� 3�7}3�ڬ`C,<2�v:�r�G<N��i\�r���<d��+@��KcA87IY+�Y��(����HO���sb�P��lm��^�*�����4�΅%�}��ȼ����`;s�5�1�h��j7^t��]9I��$�	 :U٬�9i�_O!	~X���/� � �o��5=�|(�6�|!u���tl[�ł;v�t"V ��a�8��Z
y9�	ը<�h�s�������2�m^�!��jZ:�[����!9y���[ �˭ZE�㶀ݲӹD��Sm��莇ƻ�Ë���l垧ħdׅ��i�<~�b��$�i�?���Ɇ�Gz��!�����Z�N	v5��%��/5G�|�	�]{��iW�j�Iqܣ3ETr���4���;�l�K���ݙR�Z�zn��a����m�R��5S`�P���nۑ�⼹ry-�,'�N�ӻ#����r��N����^XN�>�������-�F��`2Ot�����ڳ�	�({�,�v��Za���i�����,����:���I�6Hs��u�����d����"�xFS)QQ�ޅ�^�1����m�������?m �i$`�!�|̴��G}l/{L9f�/g��d<5L�8�@��C�����t̪���Y�X���7��ib�RƼ���R2� ��Ճ�r���TO�#�I���� 9^� )�YL|���	�2��p��XDp���@ɬ;��km�40�u#j�Q����W�z�n�L�2f蜐fu�*����x��PU��É�,�,�����K#xv�)��qӗۗ����!w��`��ID����!T��-t��:����n�����`���&^�~��^t
R�X8�f�
zh�?A����<d�9膽A'D��%��1���/������h��i�)�8P��D��C�t;6�iw ������l��A��E�6U\�џ�n�I4�4�����O�^/�z5�a"�s�1S�L���;��t\�h�g��%;@gXjf��q��PA �0U��)$@zAˊO�����:X$9l�{(t�1���;-��>Ce�����_K���v�/��w�'JI'm~sԏR7�B�}��J�N3�?�U�t��u����l�f�`���܍�i	{���ԫ�-)H��z�%z��n܄/�JN	�y��n��0PZ*�!Pw2j�݋#�Av����2�j�A��p�C���w�̟�W�;��c/6�᥵�Br��Pߕc���~����3�/qϢ"/1?ПH(b�f�#�$w@��{�ʍ�Ʃ��辶�d�� �5��#���.ǩ��Hq�w
��o���\����B��҂>�{yY}�g^5��[� ���� ����VNq�me�>�@0��r/�r����O�;�+����z&t���I7-�[iǛ��	s�g�?'���c���Ⱥw�mt�v�sL0��@�	�tV�%����,f����U����:5έ4=���%.Q�td�i��,��8|N��u�,Y�R�y�)F�����S�%\'Y���fM]��M��X���z��d�F��k��N>�䌷��������"A��R�|���nm��:�6=��Qe4�9).�\�"��P��x
�'��xO=�rf����h/�$E��En�h�U:����<�'��x3>|���w���i��3�T�������<��G쵨C8ݲʧ����I����c�ܰ,�T)�%u���X'��=�+ڼ��B�Kw�b�����`&�ѯ��kx_XZ�N��׌;~e�,qQJ^�.�|��J����vr�ݚ�k<��՚Uv��AP!GLJ�/Qh����9�S�N���$�+�XD�)�p�ix�H�V����ܦ�}H�خ;��b��\�N�#�k�M)�:�~]/w�H��������?��w,25P���Y��Y� ^���[!��vw��_�A��1�zJ46��7�~�$�ẉ�����[�����O�_f=�s{2B�kԅS�.	.u}�DdUE7���$��}�d����ú�(7�p�C�ے�@��ɧ����h���s��B)m�*�|������,��8�������l���衳�f�uy���=^@�k�_B�3齌vC�1~8�8�\ewS�T�;�SdN"���B��l|$�r>g��jc)n��tG�H�
.㨇O\��e���E$ǬJ%ϑ>A�-9ߗ8I���
}�0��3�$�T�4D�/��u#���ؔ�4�xņ�L����{ef��(�B�At�N*.�p�Ai>�tL�]s�/�o��4m�ӐV��K �����Om��ST�fwqN��K���6���m/Mŧ�]�G���7C��&�@�>��i*�ܨ��cÛ�����H��gV����� �V������+d�Z�;�v͐ǲ��ݴ*�j"���Z��mk�
�(�!�����H/IdJ2��e߂-ZLOs�A��P�%�X��`�p?W��+\ŋ���WEs��;�)�i>�Z.��BȺ��<��q�������Cܱ��V����Ѫ�M<�q^^���t)
���ɦXlxVHYEB    fa00    18a0v��o6���5�f1�3F,YГ��y��𶩎�fS�ڑ�6���%����U!��xz�l��9X��>Ãn�mE�_�����x.~ڻ�drh�a>���W��t!E�=�#�c���M\�y�UAӅ�h�!��'����m��`6����$0��S�d֝췭��,ެN1���t�ih�]��⺥H&�y�3�wS\q�
ʴ��1�I� ��~�0s$X7�٣Y��f�5���gde�T�} �f&*(1хq�`���eؙШ9P[͎���³�f1�����'�����ؼ��մ�!À�`��h',E�:D����_��u�::]uuߪ��_��t�x�#|"j攻V�di��I}���1U'�����h{aڦ��S{�!vm�:]��訇:�-���V4s�<���pMV���%���L��Jp�Duq�n�q)<U���H ��3��5�j�"���H��1�m��Q�)��[
5�(#�T�t\�-���0XYm
�@��{ۜ��:K�G�z`贏I.V��*�,ʄ�N�,?m���ͬ%�V���W�@]�@nx�Wr���SE���S�Z��p�,�o�[lʽ���d�*TIE:TF�U��F�b���s6k��6��)���bC�4��2��#����/}%�@�.|ADiݵDĪ��?F����m)I�&��w�i���u=�e�Ō�;����
G�hQ.<�i��yu|۴��W��01�����0�m���S!24U�T��r����_P|��Er�l�D#�0ˆaoY�JӝC��Xx}(���ϝ�"���RD�+��p�U��p��W�Y�C��������˳���+�����J� ��O)�[���3-�v��	�<�)�H�(u<7�*ҝc���#������"%�����gfP���O��ܒ�Y�䓖�`;���zس�sMe���H����;]��Oi���n�:�ލvx�\�d�#&k{�pr���;¼4h�d/��+�L2�u�u��T�R����f����r�������á���E��[-���.� �Q6���h⛘���[TX��Ej ��BI��+r�7:	�Qc�R�6p�f�1�~PB]r�����
�U�n�"��L��Ѿq�;�dEp
�m�3'0�׎L�_���({�^m%HZ>�ˁ�3˘'du�[3�����U��:%�l>���H� gVʹ�x������7$ǀWx� -�[I��]��I�Tw���:d��_o�g�c���eӇ��xUظ�����<���ݢ՛��5S�:�T�><������4(:�O��n�����L��τi�`-�[ �������=Ԛ�t�crN(Pe��U3��e�Q�3j����[�>g�r	�y���/��/}�UR;x�`;���9�SIdT�@	���6/�h����韓�r� ��f�6A����>�(g*���U��<?�6� �wfޤW�ds��C�����2�����mx���1��2J�h��K�������V��V��;
����M媬���L��ڂZ)j�[���<80͗`҉:i���^�ud�
�/����oN$���=LQ�θ��A,x�y{~?��w[տكT"@�b�-8oǨ�zF.0�]� *YR�+�����m�)�fa	/�s�P�GT�`9���B�?���^�e�����as���v���i��jB������S�A �R^f��3�Y����/T��M�.zA��A�y"��)�jp}��eJKJ ���{�	`q�W�i<��0�~^�Eq�@�ەI�Y���1i���4#8�&tK�:��3v(���Yx}v�ê;�uc�A�@�|��,×G����S�K�o\���&Vt�Lv��,[�Y�������6�����T�k	k��@�ؤ�þ-����%t�N\�F��sLN��3z�tm�oF��fc����[�L�A@��н����/jG��f�ߚ��ݴ�.Kԋ-��N����֤_rM��Њxt�4��jǯ�G���`j��U��;ףn�k�j�=�H�kS�դN)�k�Í�������З�ab����F�JhnlQ��q��h���;/��.b�F�#
����((���D�����l��AgG��'�Bk��6&,>�R �`��m�^�5���ȷ1�q���$sh����r��e�V0g��A$"\�SJ9��� ��-���ZX~ ���X��u������E{�۔�-�椃!^H�|��%���Z˧ɖp���f�t^�ۆ�w�|��3���8��ԡ�X!�5�R���1���@�P������RW&��x2��Ն�f}�Ŵ��/��jJ�.�ٿ�d!����ު���q!A^/�X���ͪ1��kRI�����*r��� IM^�u�N����6�^���!�o%p��JU��z6�oB(V!��ÌY�����{P�����F�R۴�7�]�8x�/PD�TF�.�`T�Y�ܔ�����B�-�U���ݱ�j�1<>�J1䃡���J�%���F��/�+HF�w��g�֢�(�[.ܑ�+���Gx��F�k��)xKej��O��/P$T�r�i|�@P�����[Ǭ��Op��u�]@=�>*�Lv��va,:��tl��UqF�;�:�`�O���%���a6 .�a>:>d�k�2�ﻺ1�C��9��mŝ�ɡh�l�������o��vp�-�'�d�d��Ԑsg���^�/[�]~���?N<��r�,�����H{�zF|�G��/���V�xӰ��َV���5跘s3�/y"�+*�]*�����o�������I.]��q~�ym���⡫���k�'��U4��Y82���v2k��-�+eL�+Vr]@HCg �G`g#rh�:	7�n����ӱ���W��G9*˽7]ު~v���9&�h�+{k���/��=f�E�$\�Êqt����������T�&h�{6%*�N�3`^�����o�j�lY�"Y)�(csAL�}�p䳁��j�Q�X=C\��cZ�v���G���P~��|�\5��fpU�Z��Ѓ�5w�+�l�H&���D�b��'�@�W��tùU	Bʾ^�@�h�iqyf�'���o����"�z�Y5h�2�KoA��r����1㏹��;���I�i2��m�'��ͺʜ��E�+���'�9�.��Ho|�>����OE�����^&�w]zk�ܴ/BΓ��H���41Wx�N\�+��|�M�w�ů�"j��m��Er��$SP��y�����b7��(��@'9ĥ�<���������g)���j���4�m�*�˘�l��j������\�7���l��%l�p��4��b�=r�K>3�ګ�8�I��k�]��Bw����@Men����|vx+�5,�z#������G/|Xq2��c6��S঱�7����ވvȘ�����Ty�A�AQPI0d���#�׎~��7�[l ��',Y+�jZ#ekIJ�ٕޞ�.^ ��ߊ�^��b�î���`i�ٳ�i�{P��jg&�׺p�k7���̱�ڿY�SSK�~ۛZ����%�u����o�L�s�G��o�:�L��!�c����l�z+}٫cuAD���rΔo��X:�L�� )��>S�	L���ri�%��;��H��U7��_����y-q�?<� |��n�:��R�
ev�:��O2sN��|�gu�a癟�֩C9k9w�ŲM��2�O�?�3kQ��أ_��H�Io���������v@���d�zZl�����W��l�[�Y�5DJ�DC�5B�������H>�:��2|n����Qs��X�K�\���sZ��(@&9�o��n�U�1j�0e4^��9.�~�֏jyܚ�����EA� ��r\I�suzbu���bɺ F6���[�Q�����6��7=�S�I�(ط��0^57+×;;�js�~��q;Y���iC�#�,mKk��7�J[��i�2x�,���8���yOr�ߍ���ZݓK�'�־��Z��W��-q�Ąh��8>� ���C`#en�4��;�D�\F�J�g�@��F>l��<:ݪ2+�/UH�!2��ж�����dpND����u�
;�EY����g����Y �K��;�����܄�TQ��AI9"���G^-��#�pn�k��Ѡ)�[Zd��4�G��j���h8d����i�%���'��������<N]�Co �@aG�.9�g���}_�>�3��3�jY�<�s \5���N��H	��1�&�� � ��ug��:��n6#��&Y������rI���7h�� �`0+�`����K���m&j��2U͐�Ik���؈6�3�9_L��{�?�@vP꺳ؗ����)GzBk��@%���Kd��.R��MSf&�fN5q�%�%���وg-}�Kì	U%;S��9r�-A�v��&%|�we�������K�辷���gus,@��P�"��.�tNE�,�e���2�)�~�`������v��Ͳi^Ƅc��)�;�1�A��j�J<��T�k�B˓�"n0I	�ɫ�0�e�{�m��bϴ��uA"j�$�j)!�җ���"����9��UQ�@�D�F0�yi�u>�
t�k� ����\<���#�ߚ��\��@���o�������@��%5U>��<s�x/Od�{Z�����[���Pڸ�6N�ZR�?〗2����	MW~��b뎈A^��2�|6�>��y~��;43}ѓ��7��a.V�v1�*]�+wT�	q*c�89�_78�[��'A`�5볂t��7�7�	.���4s�ɳ��6�o��X�?:ޛ��QJ��X_��;���@ܼ��������
Y�ʾ����V����4��q��6m��;j���"/��$ǓD�>�%�v�)4��oV4�&����Y� M!����i�Y�1��Bۍ��%+(��a@�J_o%���V�E��� ����R�	T�:KeX��~�;<6�"������TwC�X�/^�0��o���)\NNƳlܦG�,;RL��X�p���Ĭnb�d杷����i	�-�siȔn�-��,h>�4��T4F���'�9��.���D��S��$���u�n�S�]�V�ɼ^��m��ܯ��>:�di跟���{����+��@� v����V͘P��(����!E�����n�qj7��_��@�4Ci���u��{���}{]��+^�N�Ɲ3a�d�����7�v[�����){�D�j�2�&�y���B��'�0����Yy�ӯi����T҄~w��c��7s������l�U�tH	p��`nV8��~��ݨsJGfd��~'�N��z�	p���Eu#�p���� ݎ��v��"&����$�Sy3ȯ���m�f����=�X��}�i.�T�\=�{�4�4'nI��{w�Q�v�!�j_��X��aa�U�����z��7m*.�!ks�b�ɆX���J���2���EO��H0siq��٩�����5��;պ6W�گc?Rغ��r�$i�(IMG�D�s4�aFGX�/������p��3Z����{��?%��z�YH�o���ҋ�/L��C�������6���z����*��L<�������[#�=٩|/����W]��4sv
��=�e�N*oW�g���������ܽ�� ��[� Ns��YP���CB(0Fk��� @�@�S�߸\�j�V���A��6JUg&[[�ʜ����,9�� -�D��3�%z4U��@��H�"�dZ�'�n� j/ې�Nu�޻��@LE���zPq	���h�������i�j��.T��#qZ�`��T&�bKw�Sa��:]1�cb� 6v�{�\�G�+0 ��pL@�^���ټjn�a�k�%��-�*T{-��dk��|3��e\�jw)*����*���`GT�!�Z�����������nՌł|�?��f�$i3S!��/�& �RcÕ�d�����C�M�c������>�
T-��y��-}TRc�I�]��΍@�%���Vܦ��
./�!���X�T��Hʦ)5Y�����iU��i{��>Cz�?��{
*]���7e�RyY�XS�c�M�Q��L������^����+��XlxVHYEB    fa00    1200�8���#j����bkNj{��6�
��v�l�y@�3�ۨ�]Yf�
R�L��)�>8����FR��5�tC@��j
�UJ��g&�ǽQdE����O9��W�B�:i���t|$��Q���B�Wx�u3���Um�q	68K��FTn@���A�"�a�w^�`i��- ��9G�+ҟ��(��̄���P&�~Y�JzH[�[���'I���5䀊!!�Q7EM<�g��/�����Kר��/���-�h�W����B���B�"���T���{�����mEv��j�=�Ť�g�ղ���옻dW$�A~d�ߊ��S��b�!1j�7�/�m
�/�;����ğ�9�b����^�"�'�pK熶ľ����+.}<=D&�6E]�l����h��nV	�^O)��'���L'�]=?�c@��%1�dw�Xũa3��EȻ�e]�
�1��;�D1��)4�N���eX�WX�H�P��
-ԃM���.���-U��k�W�捁��m�V�ݳ�� w-���08<L����0��i��6���Z�+r�d��,(��U9j:����:��[Sv��)B��#�O�ЀŲ˖�x�G�JK���|��^�)�ə C2�]�S&�5!�V%��A�W��,qY`2����+9A#�i������Ÿ���Yy5�xw��RڋaL��������������n�����Hg�y� �d�/Et���ړ�N����b��1%�7��U��85ن6=���6�]`5�ǩ�?�������
���G5��ȹze�2�.u�ć���r��`�I8/()Sz	�<�g�І�T����V+:UX��P/�5������v�����Ǥ>6�)-c���'Ȟ�|\�%���þ�ؗ8ҀL��o�����D��`�}��$y#51Y�4��fl����)�f�_��|�����G��I�&ɠ�|�D�u?i�I��=2�X�B�/���k�,�{a����0�6���~#��h[/O�6g�u?�-�E�q���M��M�Z���*n��s�7��z�r�=�C���9��G���N���h|�>ΣWHr��JF�>��@����5�{���u7��I�h����1�6AotM�2�o���w��Qr�x�BV>�z�{OnS�ib��]gFqAH�v�e�ܑ{�n��GJ�x_�>Т��mFr�ϟ� MIJ�Sֳ���VL;0{��4�)� ���f�G�KU<��3�r��g/h�����y�6�}����b[d9�ے�ڭ��,�0����ٹJ
J�#�\#�<u��d�f5?�75oq�)���%��ޓ��4���L9s@�
j`��j���B��,�=�)�
��U�8���Q�Q���J;�UⰈ�iV�ߒ�vK���d��(�%S���32nt&��a�d(���Z��W\�_��6�k��i�H��.b<�k�>���C55z��g�A��	һ4H�rD��A���zk�?A9�����~z���$�@�+�g(8���]8O���83�n���� t��H��ի
��f7�X��pG��z���_�J:��&mt?�whaPZ0	��/4.��z3wUS�>rR��������k�;\�Z{<��y��%���$/�Y��X��?���ve���u�q�a�	˕|�K����$6S̂ڿ�:Fڑ*�5s\����^���]<�T��@I�:�}RkIų���W��se9,�yD����1��R�QIb��R����?M���7>+��0�S���OU+H�쁋`4��7���,9c"ԥ��VI9@_�֔�fdc���>��z�#ܭ�)������|�Gu�����@�V8ԕӪ�H��!�q�nh�^�l�ә���y��'�p��i�Ս�x��8ѕ(�Ss� [kX�!�[�A�yw�S�6Y-�������d��k2�;���uI���%��p�ѫ�̷�B�䈲Af���H���%��Ϗ�O�\�cp�3�p_��>F��&9���O�[���iބN�7��E��oA��s�Kr�[%��Dw����Ξ_l�ePo�U_o�7��/.NqO��/���]o���0�\�M�|�+�`� ���
2^]lj{iuw�t�}�Ⱦ�P	������r�B�G$~X���?7<�m�V�%"�9O���W�d���t�o���A���� ͝^�q���t��C���|c.e���ؗB|��S*/��ɚ YV�r��e�xE~�@i�,�����+��(�MC\�� ������F_k���Deޢ�ۘښ�:�"�s��;9����0	o�5�LT��,��f�t�i���n�Qh�m^�%J~c_��=��KJ�Hk$�zLmj �'�ZbX�s�����dK��Q�0�s&�}���
�,��9�kE�ܮPU�9�a/X�A�b7Y3��8˃YTMꓔ)=� ��=P��f�*Θ�A�x1!|K{5�A�����E��mhW�,���w� ^�~e����L�C<�x�ʽ֢���c��gQ���]�^,��!�p�aˑ����ѱQ!�tJ[���C$���N�4��w8\[����69�dF��R�0r-�&qr�&ͥ�(���x����2��]:G~ ����<뱔5z�lw3w�;^(`.�L��}�BMreh��:u�J�[�Ua0!�^L(<`�2b3�R��ڭ� �0�P���R��u�z
�HϮ��ʥ5q<�z�0���<��j�~��d5����	�2D�y�X�����땼��ǵ�7SѐD�4q����~�.���<��p$�@���Y�E�<p���L<�d�J
b�~�Z��{"��%�&n�vL�Nw�a:+6�f��	I����=���U�b��)"�Xm����掁����k62D������h�u�!ν�L�~�+r��>��������I�ñ1G!�ݘ�gL�KuF�LB\���g��!����\s��b?o:TI�{'�;�J�p՝��O@./2���W���C3���{Q�/q��{��c�MKы0b+s?�M7~�d��0qA�ϢN�SYkh��_���`P�R00���ySI~@W�0�B�V^���+?��[��:��zG(aS�����(�P8���-Q� ���=܈]�Okw�k�Z��i\���l�V�A|���f }=iR�e���;ԣ�Ą~T	a�4y��l�/Qة�iS[%�PnqE�����L��������Gf/����&-�R�}��+򾵰�� �ʥ�����;�鼶J�Yr�$�d�����Z�{�Mo's�����g�lC���ƃ�D4g������m�����}^��G��6�P�d&�;,'��t����Ѳ��e�%���4�(��LP<Q�cY6گ&
J� �D��� /]�"�����*�d�g�(":A%��iKCD�(-Y��{BtC�iL��Dq���Hiۃ���L�Zf*�T���l;a�!=�;T+݆�:���NT�v?�vl�F��Csd�M7kM��Ǵ���Bzk�R��Ns���~ƞ�r�g�,^�D��{��@0Ǖ��Y���s=����ԑƔ�h.�=l����Ϝ��3� w�x,�>���	r��dYC��c���&u�rqn�х�ڸ!A򿯶&Ah6KA��^Ž����/e/CG)ܯO��f�J�0��[�:��&��/ �����Ҫ9�5~@nVl��{����0'�A輬?+�]�-��R��T3�����.�r���2���4��3ߙ�_dZ�eB�Wأ�:��D�9�v?^�r-��z�m]g�E�1�����<��_����e1H'��(|Q�0H��}^�c `�%�2����{�P���x�>��x�.fE���]�+q6G8�����y8_j�	���l�4 ����˟�4�*�3%Ϻ����}h*��Oqy�8=(�A�_C�fr ����=V����Mdq�ط���,��z����@�����2�0�t0��r�m��N�a.����
t� �����\x�:·[��i��r����C�����'�ۜă��,XGF%��k�;q����1X�|MZ5Zv����S��������Mɠwm�3�Mw�X���w�ġ�(���S$
�����h��~�,�C���s�J�.���Ӯ��J>j23+2zZ]3������ƴ@��A*?ٳBGz��T�R�����;9��(����=���
1k��0`�h���.��E���/�Ä��&@kv�6).q���g���?L����IL�z�j�hi:��5L<!��NB��~W��R�=��䝠�C�^(�N�?�a)�ܤ�;��Vᩜ;�V�Bp������]8dKꧥ��O��_S'o$ĪW6f�[�ݮ�g"�)���+�$��n�	-�g�	�����c/�p3"�Y��k�9�F��hr��`����ʍ�i��;p'���)C�6yĆ| n7�;&�#�ZΉ7�~c�L�C�����=<A[��z�NE(�\rjnS4Ht�7�ź����I���E�O��ċf�nD��|��XlxVHYEB    88c9     8f00y�UԠ��Ź�3؟z����W	�$Y��_f�B�?�)A@�ގ2���%������c-.~�0�"�}��Ĥ�OIӰ.� ]��-�K�By��A`�<���T�i&i�t' {�Z�Kv��|J�6͂��l�5:���?�o�rsG��Rl����"xt�׏�v�=,8j��q^��?fG	�jY���)�\\�W�<�`�ՠ'���Qm5/�2����(���>�}���u��8� }2v����򡮱笌ȩ�d�ʵ��!��4����ȴ�u�)^��R��}�6�og�u#��r�C4��}�V��rz$��ܐ4�yuf�Y��"���Ia����������� �d�����RZ��\��9s<I/�zkL�S��o��m"?���w��7�y��e��Kh� �x�<� O���v.�C�܄�'�ɿ/w@r�a�SP&�/���X������� 
{-F"I�HaD4���qO���9�Q.�_����� �\k�*�Z�~	��V�2�˼mhh�Oʊ0tS	�C���%��j�R/��2�E�Dhd�^�(h�p1�=�W���z�G:�ݩ��	�rN�F1j�;5Ņ*4�A����x�6��$#��H�?�m���& p��c�x�n'֪n��$�����N�iX:������C��%-�v����/�.ԯy
�
9���q�j�. R0��nZ��^լ�B��]����ȉQ��ks�GK��K+;�&�Jr�cu�I���zW�R_�,+{����G%�D�2O���h�P���v���'Y R��X%��eA���j�)K���L*�G�Nɕ��"�2�{���;A����V{Kא�1���U��R� `�����J"+�4w���)�̻>�w!�r�����J�.~g�1X�u���Iv��� g�A��Ok�GN+�5�1�L�@�"f�'C�Z�_�dr&?�1c���iC��0:	��c�2 ��g	Z�$�⪷�@?�<��e{��(+�Z�}1(y�S[�6d�se8�@4=Zu�����I��Y�G�l�4�7c����m/Q��I뾛��8\l%��8�r�>i� ����U�br=b�m�r�}]1Ϯ#�^|v}�J�8�$�W�W*ǔ���8ǎP4I�X�a�1���p��Ϣ��[��ZL^�%g׆k���|v3���w�G�b>!ύ�5��:�Oҩ�h���C|yXE��������1������3��]w�.�eez��҂׈��0S��NsDH�ʂ�j5{9���%�5� 7��uJ�rlG)w�pDWc��`�U�U�x� qV���>�U��ecvӦխ�btޖ?��࠱�����!lw�0�'�t�q4���Ky�)�v�5㮅��]��� ����Ac���#9��+ce5 û�����=�`y�*0��)$�w9�|��GD�wO���m��bUi�b�+/w�.b[�MK�Њ9����cw�7N��8RC��j�hG�c=ԙ�b���U�|���!��h��z߷����W7wRI�@�?ߌ�)Cc?>�@��dIja�I� e��:f#�9����z���k>���*���R�.i8���-g��$<��/(�"H]h�I����o����U��ih;p1�7�ō��	\�U̺�Z�� z�9ݲ����m��})p�_�QB^����'���@������;"T�~���3u�bN�Ш��ƽCyW\!�}�=d��R������ ��6ɸ'h��ћ��Q]Oȍ�D+� 9�3Bb�5Y���-w�\��X�@S}��\�3s[����$��"���,�����^6w�. ��b�.�%L�),B��*՜c������t�L��>�$θ��`( ^c�$�--�����*1��l1����Ey�E��*G�����$�%�K�L>�CC�#i��Fް�Yԛ65����N�:�0``��;6�	
D���k���sY&S
RU%W����dZLj�Ԥ����0,!��<'Qf\F
xÆ���紴>N�ɚ�5�&a-@gU�U.a���M�/�]aW���%�ޕ�H��O�V?�xw!�wsDc�ZZ�>#,����@:�� p!�e��^��A����K;�	Ǽx���f�F#�B���ӧ��v�����9��}7�yq"��4�8�G$����|@Ɵj�6����Ut��A�$bT�9�C���N3�	�A	4h��Y%+�_ cgm`R9��