XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����RR�oY��y$w辡
"��+m������by�¡JE�.��x�����ɿ��L��[��Ws�]	��	4���;����@E�\:�۲%[0H�����"��YV�V�1�SD�ٛ��l�`����Tھ���[�Az�Bj��涶�w����;�,n�Ȗ��&ux�/�����u�E+���2��fA
$����U�����I���]և�z�n���19!���
�2����*���HA���2���֔��0�1��:�vP�_�#�~1ǎ��*2D��D�MkV�5���]*����̹��?�#gzmO�.�s���BP��bԁGœK"S�\��(��L�����&oH��3~�}��o��ۀ?�DS��R�1Ne$�|�D���
��>��3�e�&�љZ�9ڈ��u���#<�p���d9�3�8R���u�;�z,�=�fG��C���&�ܬ�V��<�tT�m�
d����eE�/B��X�(֓DB6F#�Uɘ4|ݸ(\z%A�-��"<��{�\��\0b�pL9���Q�x�8��0$��s��QW0�r8P�������y��.1�AI�a����o��C�M+��2�Q>��`s8�TGv] ��I0y�!N4j�Y�h�q>�E�O��/���p�\��N��)��tV9���T� �i�ɍ��S��72lF��>B:�$E2£��1���"X�#L�?�&�kA6���X!S�6���t������gѳֳXlxVHYEB    4089     e40�=� ͽ�_��:�w։E_�' ;� Э �X�)ȭ�0`��	S�9���w� Mu�#�� Y�Y/,vՖyqZ���l�z[+����q�*�\̯��]�l'Rl�(��v>��PԾ�3�Iᧀ����-V�0������JE�-��aM��x��m����y��؊ �]�!X������;��J��{�G-0;�Pk��ן�,��w�Ox&��lEp��O�M�+�{.��:%�.�1�h��{�e�n��^�x�=�,�#GEx��Ynέ����7���ZoS�=X�e�����O�T$��o����U���Y�l�M����ad�+�R�~c��ە	���y7٢R�-�j�� �,�J%�	#N,��X��ڥ��r?M�#���`��Q�/~�ħ4&8ibm#�4�"<ė^���D�����z̨����n�������u���S՞x�Pt�Z!$�B���7�%�n��Q���G���E~���V�x,�t��)R�5O��hD�uH>Y&�j!r�@d���\�"ģP����Q5�x:�o;[J�Pn_�`o�P2�sf80L�L�,徨F��=6.�������M����Gݬ��K��m�����ؒ����{Wj^�h}�+o|?yZ�>~��axE�9������f,�8�qnX���F'��Pf�۞�榯dp?������0���B�_��b��`0o��K���â�.?:(
��K{��j�8�g	i\�@䄉+��~����O�ߴ�k�J��#o�7${K?>�0&)�D����H_�����Y��3�Ec[��*Z�5���:�x)y�o����0L�-��Wh:��' ����ҋ`��%�dE<O�Qz�Y,y2�M,w��B\!
�b�̾]���B_���@E��"X�KU��Rd��x���QE>��<�-��G;�9%������/��UR�YKiٙ����=��d�ϏF���l���@_'DH�h��J�a�T\�}5G����W�1]�=�M��&���-HMj}� N{�*�q��YѠ��P��
ٹ��-V��=yS٫ۯ�o�6�]�:~UL&�_�I��0r�ҥ�KY�(��p�R\����i�ݹˤB���i�@�]����f&�mw+���F3�AIҞ��ukr�\~�胝A�ŵ�&�7"�;&U_��q/�U�6.��Z���:;�����(��D#s�"�I������ؘ�#���0�}RR^7�v(�O�����-'���R\W�;,�A��������6�5�D��<e|� /j����NY�	��.� նv�$IM��YۚKk�>\��W��R{\��6C��4��\�z�`F9�
U�7��j(�H �$��[��j��rNS�jQ(���>�~�����#�r}ȗe�P�|����jd'30����r����(K�X6q���h����Kk�k��׍�u*��7�چZV%#f�����	�QP7���W(�I�P�v������%=Y�����YGM=�������]�=�\��!bv�����<L�^�=���.�c���{�q��hB��~t���5:Hˮ�R�ށQ7�j`d:�4.���@�/���u�����T�z��s���T?w'�c�.ۘC���*/
�N�x�9usN��/t}�O�n��"tE.��������h>J�����JNy�5����ہt�IXa��r�P�b5x����Zh���3]�B���
EW����"�IK�FE"P���ޚ(˒i�m���1����E`Sذ����)$S׵���0��l�:� `��*sw�RS�}��Ʋ�F��|��bR����S�d�+$��u49��F�y�ZF���sV˨0A�r��/�~K*�3uD���{[H��s�R���7r���n�' �� V���/t���
��!��O�Mr�T��<��?�P���E_R�4���Ť>�0hfH��^����A��~�h0�G�s����"�T�f�ʝ��AC�ք �}\�|HQ�R���Wקʈ��鞄��)��8.{A��S3�H����>O�����H�̮[���x�x��4��;�+�g��ĉ�xFU�|��i�Ͽ�"����F� G�C���S�lup��Io��z��
��q�ƔNr{�n&G�m�l�����{o��Wu}8'��l.0c>x���'k@�1ui<�Q�'���q�.�����v��?r��qP}{1�XSm�J{����[�	�O6��>ϡ��S���3�Cg�W휒 >+'k�� &�V�T#�9�Ѷ��ע�������>z�ܼ��l�����Ԓ��q2

#/�P�`�\���7�_3´/����c�T������%IyӥJC%��|vP/y��#�k|�9^8�b���MA��a�� ?��{Ly5oy���O33f�(�R"�(���"T��~����-������K�֬���! ͙�2%d��!¼��@��S����J��z�X�|J��p�����	�|#����-�/��s4��>��D���&u��X6�F��Gbzx�tDT���Y�^Q���	�{��ן�e'�P���C���p����Gy"�jt��v�1v^�N4�D��-�N��]�}����/���i�lp����e��IR��yӮ�ʁmRW��"�,	�S�4e���¨�KX��@Ur򓣀�bHh�����;l$�5˙��o�ך�Wq+����tiV�������%\I���ߐmn�H�{����p��/�����:c��
�2"0��$��+1�"�������{�op�s!e:Zh�!�M��w��"�$�qE��#��d%X�_���Rd�*�d�*�`�_��3p��Xt � �(��M��b�\f���+���X���TdFILba�����u9�+�G.S~v`���{Ω�5�<\�5�<�hӉ�5�f�Y	R$�ʷ���ʶrD ������W�^���w��^�,4k4���Wc\YMx�����3l�Pf�H�$r1�]�
`���#i8k�?: 7��-��S�&�x�=�����L:����<<�DE���ѷk��T�����#7U=ɿ*�Bxi��U����L���'�i�;Q׋�{TP)�!W��� ������x8�=
�,�O�f�7�����s�������[$-�<'��m�/�3�\S,
��-6�(&���fT�i�ʆ�O�F���(���(+�B�K�q;S�e�'q#H3���
+�V�&�	��ƃ�袘V�lG�>����ַ��.���>�����W�,�~J�5м����3}>`~+��PA�b�Xµw��R�ܤ��0Q�V��'�a��w}�@�*��j(�����U-���#�k�D�$�;�\0iÅ�_A¸��"t]�!X�o�^�ܙ�ZR��B����`��$�5։Y؉{�dN��2ਮx1R�-���l���?03���pB��d����'�1.X��U6Y>{�啪�j�cbÂ�1T���X,0/�:��а�{�`��Nіގ���X�s��S����g�8��f��=����r�p8O_����i1�2ju3�3[+��4r�x?��:o