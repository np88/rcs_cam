XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���B�کy���bQc�*��њ.g���YZf�a"�a�ʶΖ�Q��^=o��G�Q��[���@��':�z�P@<٢>ѱ̹�<'�~�G���Y�F��G�a4cP$@8&�vJ�,�����)1�
@d�T�s���
1�n]�?k]PR@�l�yl��ͫ�em�"	�U�b�lX���אeޑ��8fɬ �Y#ϻS��[]g���K�ӵ����n�nɉ�7�ê����z����=Vl������7]%�Ԉj�q���b)7��ꋂ�8���t����9O-([�����:Y��'�x�l�2}�8Lh��dw�J� �f�.�jI��M�*Є8��YP{sP Ɗ�@��]��d��;�M�*��佡X�S[?=�����B�z_������-�����3��F�F_
�j2oʡR%Po24�DFM��(@����������h�W����8��JdZ���&�(I��`��V�҃��H�'S�@H�����o)z�u�Ch\|���J�v�bw{G�7_��h���ѥ|jt|{3�<�g#�Y���a
m�N6k:,�~�;��Q�P�v��3��D��_���@��i{��@�׳��)�2���OF[<u����������::�&�j��f)o�����rT�zNÌ��d$A�!fl�����۷6&37����Wl�@L������K5d���(�L�����Gc��_�M��I��Zq.�����n�i��t�{�W������"��z�=�����m��XlxVHYEB    4fdd    1090\)�E#�%��<F1_/���J_�9����@
�r�r-����B�.�c��
��%T�2�Y��t)�v��f��Zu�A3ߘ}��N57�΀}���Vq����~f�2�Og�����v�?�V�1) ��.*��g@/�hhL&�W�Ǳ�]�郜����}>��G`�)�{���$L��eV�H7��L{ܔfQ	�פ�?:�x�%���KUe/
� �i��4�$���t��1���滰��H@x�҈:󼧞Q��=#�e���>H1X�˅C䵎�䶮�Q#�u�Q���k�V'=#�?��^�i���3lG�ݹW���B*Eڷ�����R�I;��{-IO6f4���|OZ$BF�zG�4�r�$�l(����o�sYN䠸9�Wg� �W��5n't�6�LGH@�
��7E��/S���o����g�ͲS���Ruh(��%�L��^h~��l�mnu٨�$s�f�(����;N1��#Uk��^�g:����tC���"|˰���qh>p��X'ِ}Q/��w���:�7f�W�0
��3#3b��_2�VZ\3-��I�����]vE���H\�{j:����	�5F��m4�s6P���I�8�9
��Sg�������	�R/��W���9��W
��#	T�D�F4F;NzS�h~�l@����~&�m:R�D+���%�2bM	�7���?6Vߏc����g?w_�y��Cѳ�����i���k��:��X"�x�������:jv�:��|1�i��VT*��媟�F%��<��Z7]�^X�G9o����ȁd:i���횓^�w@���>���)�^�*�b^������s�ʀ���mi��z�ֳR[<���tBq�)�����^E��"6;�Fēн��&@/-��9aw�<�Q류��v�e+��!�>��xL��6�Q7H�=�t�zg���wUD��$���0�Y�RkV��T���e�ڟD�;Üs�- a��F��Xp'�6�m����u�����Q�L��|�=�^j��.�,N���C:U�"jv^�	�d7�wLc7\��$,�.�>��8����`�cM9 �� �PC�E��.f�蛪��mxJ����%'<$��R�4���=�݈�z*�J8�����N���6��S�Ξ��D$�Zdn1H��q&c������ky��_��mkk�V��㺒�w�P�F-�΄� �� ٠(aȦ"$�4W lJ~ �� &s������)�d�5*�����ܶ�?��Ҙ�+�/�&����<������-��-�e�Qv�Q���,�D�qy������OR:�-�A )���=�� ������y�d�<����6N��
�AFR����[\�x�ɏ6ơ�Z�sQ
�@6�D]���dqsL8��>�ZNۭ�H?�Bs������E�F�CH:$�Le(avu,v��O�G<k
�;C�ݚwᨻ�����}\'���˙'z*Q�QT���͓���ώ!<��v;�U�%&5:,��Ψ��>!�)�;�,�8� ��2��=�Ds[ﵸ��lR�wcJ_����{ٖ��C�B��P�(��NU�0�O�+~k�Qu��+-�.�o`����E��o4n���2 Q�@��G��:���A=�5H�,z"�d��s��o���ӏЖ��(j��l\�Y-�*F����?)��B�{��(�lW��--N��hL�Ǽ[l*�<�N�i?�
1�v��
�	�Y�	�N�@���y����u,;��l�U7��d��Zp=�>WZB`��(��/s��ʭi]S�P�Ԗ%כi� p�n���R��s E����x�)��\�f�}-E�(�b)[��R,2�.\ґO�L�V��k������ ��~.����	i��xl�&%�R&!n~E]Y)�Ro47�o�u�)/��������I3g~P�$ ���2�{C�3)8�)3�����o���Qv�J20'�D�( ��˾\^��[U��.�nC�.�!q���aG-��ˉo��|������l�E��ɢ�(�܊C)�V�Vq`c|�9�6�q���ɮ���t7�pW:'f ��V����v��9��s�[W�R?\k�/k�iS'������8�F%hƎ��'WqQ��?�s�����E��G�x���%L7��ٱ�.�%���h*t�т-��G��7}L�'��i:�����]}J�34�'}L��P|w���)�רs2u�@"���hFaV~�7,�_�l�'Tܜ�
-��.��u�G��q���bCR9,E�w�� 'ϟ�����*��]�s)���.	:�"ёS`>��}b�o�J+ҁ� a��5ZΌي�;Cty�F*���Ɠ�2�C����,<����m���^�/�������\]��{ h��x�hlH��N%�s��%�������#z�A�j���;������1�G�������x�H��x�E9�����僰ۤ�09�%w	�;��Xu������-��fC�3�(.�>�� ����%�� Zږ0+��1�+��y vD�mu�����lx�዗-Լ���Đ��8x�&�{<�9��D�l���<@u����K8���b����އO�0��0q���FM��sT�P'A<�厛�55o���^~"IN�۸%��g��X|���z�t\��D���Y:��n�����0z:�j�/m&�KY.M�e݋�|�[�3���b�K�{Xp��cc ����c7�~4ז�pF
��w�G_x!�/;��_B4K�O��cl:{+h�5��-��X~��;��,�����D���	��1����(i�b��j�[�i8���!1��X�$�#Vu��P�kM	Bp����v�l�-���˙5�~����x\؀�$W��	m��o�qOu򍮽]�
�i�V�V�f���'�vOHR$:$m��L�-����n�NM���ϭ����W�z)�ֿ�<��<(�x�C'����������{�N�+wj��`�zǲ+�H�s�F`ܝ�G���Q��`�ٙ{d1���%E���u��p"�F�bb��[��f��N4\8�C6HEGID����`|��0���Y���"[w�;��-���괭3��`�^���L�րH�	�.>��qf����渚ېʝ��r,VՃ�WI�N��@�s�E��8��U �MD�Fo���+՜�E��i��n]x���%���d~�X��g���P��O��`���v�*l���aY�h�����7����2���y1�>�?���B�r�mV��� M��֚��������ϳ�!L�E-���qG�Ӓ��A�y�{*[�W����πΤoK���}� �:�w�9����ܩ �>:,��{C:!0�#��WR
��3k�H��2��:����@T1�_�-6�~Q��RѱbUV+��G�覩A���)F����ѣ̷倥��O��4���Q�b���:S/U�A�޽'(�t���d�b2Ag}�Q��Ӆ�������nr���eS���� \�T���H��#f��5������O&��Y�;E�O��s�����0F�+���tU�������1�����P/{!w��A�%R�!!ղ�|��/yC$����3W��#O5�\H~Ѫ����L�
�kx�6�_Y��$�dn��C����W��)U����&�zΙ����>0���<���H�����S��+��%���(b��2b+g�-����X�0Q�üAh͝�jyuX��E��R�q����E�_�����#���=/��_�i�o��[>;���d#�e�*�0�v�	���#TyFh�&~y�o��W|�O�͹��{�>��蚘�.h���+b܎�OO�>��@n��P�J�s���ΏR�Z �Z���eb	a<������6yx�U6�">��d�!��n�-���J�eYN���^�0)��t>���m�A��KK����/$��*O��
��ƭ.s�咩9��
SV��R�������i|$Ux��m\�ċ	��_w|mA�7�|�J��ɓ��,>����a�����9���
廇�E&��w��>�M�\S�B�2X� �Џ�03�������fv	x[�D2+`QZ�X�攌	4�xu��ݩT? �Ho��� 8�)��}����6E� ��Jb�Y[XhG�츚�_�Y�y�(�p�C�G��