XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��[��U�0��PG�Ã�A���I�B�dOKj�	�xrw
Jv�6N{6Z���M�pP3��uI����.ią��`��:���V��S;i���#�7�P�\�M�l�����:�Y��[�3���Y���2�q|ى�Ǩy���m+��� >�ܐW�fv��	�i��]�w&���b���r�bV�[��q�*ӫV8mfMEG����[��O��\'�L�jo�4b��<���T:� ����
4�|���xx
-�f|�v�*ڜZQ�\L��B/��ێj��G%~	h B����1���� �un'�`��_� �4���6*	3�N����Ƈ=!$���{��/E�DM����bk|���f*�J�R����g���d�Y��������ccZ���BU'��LM6�xR�`z���#5��ﯿ�!n@<v�/d����:�D�lU�mD���J�"i��I=�.�(�l�B-�El}�8!˰�ö Z�H�Ĭ/�eYREj:o`G��RzD�r��q��:����D��c7~�T[ab��x3�h���͍y�o����A�Zn��9$�U9�u�4�a@C��鵽(A��N�dl�.v=�`|,Մ�G������\n�<+�'�Q6;ؼ_�C������i���}B�3���Û5���ȯˡ��ٙ��J#a�'�5@#Ug�1�z8�]���,���uzR�ܑ[5S���w�)s���-�K���F�8{���C�P}5�;ˤ$� ~�����4x��"_�q`�XlxVHYEB    38e2     fb0�aYe���a^O�h�w�2@��3i���ƽf	5څ�����(�r _��̽�	�ѱ6���WXQ���|;Gi��Uy�TA�S�R�'�cI3Β%p��{�������[[����Wѵ�s�g60���� R���9;�n�A����qQ`�S:�-��A7��j^Xw�`�ƫ��ҫ�+�m!�����&H�����9(B����4b��&�2�w1,H�����Z���3��������n4�a���tR�u,�����'�9sP�]g,A{*�G����S����8�#�㭼��VFRn(:�N;^( lz�6wQ�X�c	6��}���Wr5	�,�G�oJ�FH9�3rB��ph^��y}R�H/Zq�X.�5�T�MB@t�v?Z���9����ݳ^wO;l0�_���vݧwc���t��͂�^7��b�\6��v���"VCmSp�o�:���=y�?^%��V����(����XY�OA�R��{�ScsE2�0�������66�T	�q�� ���- �2�Ϣl4$A� ��ʱ/o������Q�%��`��"�D��CB�g��2O\:P�R��3i\�Ä�W���_��ët<��\n��Ś��hx����įh��{�+`5ܥ�mA�P�U��(7���I�+��v�J'`11Mm�ӭ޹v�a->OzO|���H�⺦�R5w�,��W���I�u͝��ɰӄ���b�y�K	�WkܤH��o��3{ܧÉ���'�S��"rY3�{l˃/w��G$�]#���%JF�R�8���m��K����.7 ���[�j|��y3��.�O���ܒ����F	�z;��2r�H%����{��^A�(����
c�謘H�6�|T��"�k�"�5�e�Ǝ�n0�دڝT�T&F)`��_Z��y��$Q����>�u�Y������:�)�ڱj�BQ)�iD�4ʈ��q��r��S�%�%�Y�G��V����^��G���
�-�=U��a�튍��*^E{ެk�;>>!%T_���z�`3���ɯu��,�!}��!CLY�LW%�ASDq��f�W9��:Z^
6�Z@S��l�p��4������:);�_�U�i߽V��4����� �X�T�A,��aa_[ Q�����
FA(�&�I�*<E��P�٫� ��,|�a,5 / �KyJ�WdZ4|����kL�v�,�q�J����B� fup�.瑂�۩�m��ѷ��W�}WX)~�gb��^���w�u�nݩ�(p���~6�P�^��4�k���D/���k)o�&5P6�H��g�3���n����m���3I�J��\�+R��U��g���Idq����.CČ��������t�������UH��p�B���-�H��^�AZ�͏���'�m��O`�s��k1�1V���d�j��_�����B!������up�p��DZ�?$�&L��#ƜH��t��#���5�_�P�m�Yd8e���m*z��	˷e����/�c���<���dD���_��w��Ȃ�*	��� [�r�Ӄ�_��<���� ��ZN-7b�b��M7M`0����T�[gߵ#��\�W�r��v�a��Eϐ��v=,l'�?;�KƉIب��{pXN&c�b���([������5���O�=Z��id���ԡ�*��V@���m�����	H��x�p�{Lv�]�z��CZ�q�Y;��n�nɲT+Z?�����g.�VO����m��d�3Ӡ��� ō�0�`�&�+4�U�W�Y�2�0w\F�茄}A��9�&��QwJ���+��|��E%d�GIS��%sY�u59��_��/�����)�mrx���#��ս%zD�$�>�_�I�~	�J�G����J{\�R�ng�%f�[j�r����!��wh���ù����c^�e��l�rS}�XDG�Ě��b�A"��Z4����� �1N�CѡQ�Y+q�|��NJE�$���)�X�.����Q4z�)��!"�^E�%|�(U���~v�O���	b?���SClj�'�����{�j�I$Ue�[n(H�C�c�f�ι��1����^���Zi-�(h�_��Ѯ�Iٝz��lVG����'���k��z�\|�;p��>�ؚF�!4���k�B�\u��R0wHE(X�� �����F�Ap�SІN���N�U���	>S�6�����]���LPj�S,7�l�u��2փ�@�<G)��b8O�Ui2��b{�L�����n�P�p��s$�^��x�!����[0�J��R�{��@�]F����`��F���چ��M"]c'6���G^���h������J�s%X)f���5ݯ�C�ޜ/i �5�/)�8�|��E�@�=s�0TSz3H Mp����[0��0�d[��)�Q���6�{����^>	�{x�-�y;��M ���֎X��`��"�-�mTS.��n�$.�;�:m���d�Q��A8&���G@����+��#�70	6���/~�Hw,h�p��I�cJ{�mv�{4u q�؂��kb�Omԡ�f������m�Po{Ǝ��ݿY&Js��U���>C�ʲ�|�!��W+MF Ȱ#2`ۭ}w�2j�M��T5��1��߀k���̔U(	��p������l�w�S��p��9��"�Es�F��O�Ĕ_brO�Nn"b"X�#9�Q�jDI��)��Ւ����@�F�c�Xh>�4d�o2�e@f��g8e*�S{e��az�k~�1�U0��,�V���(o���\��]�����M��d:�%քk�Rm1�*]9	r3=E�m�v�E-SU��H&��Q��W� 1z\��h�DUrY�2��)=�̞2�ۧOޅ�'shd�͈��Ǻ���>���8CqV��gqi�|Ř �˳j�a��: �E2szx&�t8����a�}�����i�Y}��Ѱ����2)����Þg�������e�� Щ�ÁH�j��9W�-w�*�I�b��������N{�i'frdR���9S��+�\`'�I՘�c;����9�ֳ��^��{����f+M��͂��[Y:<�j�~)<��U��|�L�qm���@P��ٓ�w�����2�"����>3�.t�O���x�����o��� �Y?�9�ĆL����d�S4ZO���������M�d^f�t�c�5��h,�VR��)�rpyRs��Е��� U�<�a���!q1U>qu�=��`�H8����c�;uW3�*ъo�磬7�yݱ�g�ʌᶻG=�6=���_�54�~��P�P%ϑ���xC+5�B�t����������c�|�M��q����g�\?�Ӵ�j�
���ŨEE���I�>��8JTB�7���NT���goT>0sʪM$�mD��ux�\[>p}���nUa}mW�����\rY����/]����X��
cIF \����� ������dy���ۿB�W���^e�
K.�N�d�t����~>�'��[�����y;H�3s-R�V�H'�!�t2���k5��+���X�x.pw�+�=�FQ샹-��=�(>��t	���fCb�.����?%��>"��@�R��g���;VJܟ��>]B~��kh n�����t08�|:�0ad���{�v�|;ͬ��ᱠ��ZOw�$�vAQn�?����Sl"/;õ�����!�<<B�v/�y#�q���E:�����x�]��.f�̘\�'�,�U�A,�A��'��,��Y�e�:�{�:��Y��%�-F�+}��Ex�+~S��ϊ�r��qGz�،�$i�s2��"3A;,��ly�5�-}E�b��/��z����̭�3]+%ԕ0���z�b����.f'm	�'#��q�43���>���g���X��ѓ�*0?Z�l�>/Q{��X��3�`�V	���� �o�+p����J�.��