XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��r�#?�:u'�-�_���
p��]��
?�,	lr�B��ɂ�=0ࡠ)S�0�_�ثԔ�E=p؊����������E
Ϸ��� �&L�L�9�Jw�-�km[:
�����k�g]j%P`d�L��U��|-YY�<�^�z�����듴�۞;^���j��NC����2�:�V���x7�Y,��z�r�	WV�*2�ET)ج�]�Ɓ ߵ�g����l�l�:��޼���S8RFCھl��y|D�X�I�\6�;�Ѥ&�.Β��s�k�;�f4!}
��7<ߚ�<w(�?���;����FJGީB�h�ʮ$�+6�R4�<4*]��A������k���.>�����)��Z����':��Њ�c����(�n�/���� �<6,@�M���9�Hk������"���j�wQ�8�ٛ�r�V/���8�p9��g��4{*�����;�f�>%��`H�
����]�=K�;��Ec|��Pc��c:J<#qf��r���/3��!��/S�㫈��	��YU�<�\����}KdKk>OL�����W��ᴎG^�:0��8E?)�M�����_��V��ݰ2@ߵ;������r���@����H��;����JԺ�+O��8s�c(��<C�ѿ*(p�4�}8�1�#3�k��#����_�C��ϲ��O%���ý�-.7;�2�ֹ�&�\�ٲ��3�O�Y��1q)��e6r�$�bl��t�as�*�;����!zXlxVHYEB    fa00    2900����iW+����7I|��^eQ�D}7f�w�ryU�pc���w��~gKXLԇ��\�<8�1��q��0������� ���^[���x��(XCx��4�wq�.)ż?��|p�|TYrXN�0J��6�c6S�>/a㧼Fx��`�+�#u�[�Ns\b�+ԇ����Վ؎�yu3l6�7%�3L��	[�^p#&U�(�T�<$(L�5�k���}�w�	�
1e𢘺t[0�8f|��?�P�KmX���=ɗ 9���k=�p{>�_�Oj��n���6!�S�ʚ-��S�v^��R�|�>l�N�$ <��摽����#�/v��U���qWRs2�sR�w�f>u��w<X�&mp�C����懹z��/�Af�V�ђ (�"��6�h����gH��-�,Q���k
C��^2���x���W�N¬=/;w6���M�l>TE�4������ɼ �yK���/�l
�y�S�N�����1g���Y�V #� σ}A9���O�ؑ��r��Ku��蕍
x3���9*��KS�v��ᱥuP5�dna㤖A��q�vٳ41͌c�?A���Q!�8���A��б�sK{�u��h6�z����ʉ���G��-����E�!����q�͈{�{�xa���&���3o�<C����d��>�`e�˃��P	q��+��˔���b�d��纼�[yg�n]�Iᵽ��:�V��ܛ�v�9<�щ:q`^�P{S��� $VB��Q�n$ƨ�u�b�yS.�:1�`���7E)�g� ʎ+б������7���'���JC{@��D�赵w��yb�JI�,S���d03����j~oP�-�J�"c�jЖLɲ�r�C�Ԛ�EG��t�1(OْG�9GL���^��tM��3ӥ*����1����Tez��w���Oz�Z=���x>�X�x]�Փ��s��ԩ��ЗV�8#|V+�� ���
�P(�.o~)�\�Er��u�ʝ*R�Zp���#��uS�4��Q�I�asVU"Z���m�a�1��Dۘ��xr3��.�J�ө`����}�|"Ϣ�q�
7��*����+,OeC(%.Q篴[�͈�r�QU_�M����`���!|�s�(�xP_���.V*���MN��ʇ,��o3��;�2e���Lr��O[������� Y,c��흀B!�g��a^�`�3�/������`���L}:f~�<��e۽����K��~�cS!��6��J3��ZFc/�cFA���Zqz^L+���#��R޺p�OL;{�1`��Y�ޢ�gnd��E�C�Ԭp} 
��/|O�C�+'7�;��#m݌z�1t�bǙ�:�- 塠�%�t5Ykb���*''<"�LE?�&[��Nr�V�*�	"9㌗�92�Y���|�_Zęg��ѐ��M�!�Z_��q`Q`���-c͇��}�j�Ո?�?�i4��-�m/V^AEy�+�+���o�.γ�-fߤ��2��V �ĥ9�����i�x��߽2�����q�v�Z��������"M�ü��'Z��Ļ�����5��Xu�p��٣��]�L݃P�'l^�vwx^�
��Чr{��1�x� �P����#�j6%�z/�2Qx��{5kC��J�gٜq������u4��Z��O�gՉ$w�}��54�j�E�v{+8#d�,˝�3�Z��җ
.K�R<�́/��5=�:�u4��{tG��16Y~�!4���E�"�o�+�Zt��l�_���F�@˛q��� �"+,I�A�u���� 7�����
�Ƕ�&�W���e�O��Ne�#H����b6M�X]�}~�L?ky�H���dkIz�Aj�N��ac���(�Z%�U���9]�FG.0�$��8E��n #��|���!$~$�ھ8�v���}s��L���#W�N6�B�؇06^ �_�BS�q���xF�p!nn�� &B�����>f~�Q}`�� ��3¨��7����X�	K�Wk�]p��,�37��_;;N���ySo�PV��g�h��)A:�c��4�a�с)�Q�1WӔ��K�}�
Xš�K9^����z�d��ӎ�=���UԀ�;�a��,BͿ�r)�
�\}�P��c�4���f2#e�)�24(Ī�k��[ѥ�Ϳ/�OR��\�224a�9���	[ޏSɰ�phB�	���]���b>^�U6�y�Ӭ�w�Ξ��O`������["��ky��iqH���
�3�o>5���%��>j��:Ž?8V�{���6���v�3����$x\��~�#��d��6A�!�+u��[Km&9o��ݠv2�$�1�2�n����6F[�NyX״�rS�������-IVh8�~�[����2�+�d���qo������$m�4$d���_@���煏�nO� �a�? ߶M������XF?�1����HHd�AL]b�]\_Vu�5�)TW7��g��f�0�a�%���x��p�� t<�瑖�#1��S!ζ�)a�����_��វt<k_�8O$�(�Tt��..�R�;�zJ�!k�.���%_����ɾ?��=
	N�fkם�|�x�"U���&�1s��([5�.���L���
�3��?�R�鳆������ �{3T�^Eh�}����+��d��$I����%]0�<��Ij����]������hI\��"�.?D�J��/*�JCt��R���|�VJ�ZǂG�ֽιe�EzU~�x����f�x@V��՟�O&1�<*��Mª�Ѓ��59��c���S��h�a���% �}�ڕr��e/\�J�2.��j@A�����NB΀��bAY>�f����E	AږecC5��A�T�{��0$�M*��C�uҌ�j�	�Y�M����N����{�4t�(�C�P�:w���"���^s.R�ԸƋ���1�(?sij�[����E�m�Ux�������Nw)�a)�e�����Ʀ����w��\��D&�����J(48So\$<}�
P> |bZڨs8e��p4�k���*�
$����'��(����p;"*rd���~JHB��5�%������l��U��J"��c�"Fw� ��ޜl �=��*>�s,Dw.�g
�J��M�������×�����c�qk��J*�~��6�����I3�Ƹ�-NLe���S� ��6�*����"gK�qü��c�}M,�^����B{�;��=�g͗G7���:2i�� Aa/����k�/�~
d�A�B�w��4�E�8"��/�&bՖԄ����oRs��p�RSU���!�t���{�F��D���
Y��̚k7Ĵ'Ĥ��Z5�����O0;Dn�F�lrnI���2aN���p����[��-�UQ_%!�.�d�)A������~���%b�C�}��w�����M`����C�u?�S��ԥ�5���刚c<�p;�̟~��m����ݰ?���L�a;��l��I�i�HAb���^��z�J��0�,��J�0<��0u5q� ���E� ��1��m6���8,*:�q��{��_"NB}��֟[l������e�O�h���x����r��WF>T���._V�	�_	�|�|�pk�?���q�׬�jGlI�y:Tq��L��X���&^�WPp�j]��r�b[h;�P6'�8ֱ��@�):!]	���<�]�?ˮ��n�1�"z�:�K 7�a��v9Nӵӊài�l���ɪ�Ya\���U��<1����eK��̵�R��ɷ����{S�y��Or���.T������ˋ��;�Y<��T
�Ls���!�O��~{�,�W�4�@>�␲+�cY����b�R����4�;��w�U+�I|�D��/��l8�-��eęy�������!5����	���5�N��؀0�՞\5Ơޘ�dG1�e�)0�KS�S7�'�4�Y(!؝}�C�/94��>!�j��{>#�e󥾏п��ok�C���ԙa�y���Ԥ��U�������?=߮�5dǏ�~ ?�YՄ!P��!�6��=����V�������G�t�m�i�j����.+f�~d>Ygi�"���kŠu���H�"JF䕔ou���O��t�1SEy��_ޫ�� 
q#l��4�����dw����U���p��!�9�,��{ |�4��B���~��o�<�ퟤ"Xץ��8Fgp5�IH3:3b��s�̓���w��t[�V湑vM��DwYl�K]�m�F{m�=C�C윲�ӅV�����i��\�	Y��l��w���2�	�WT���B�u��A�/��hDP����Sڏȶ�m�_��C�B��3�{s=��!�ӯ.�+�5�D�8���V������O������r�o�.hr^�ݩ
�o�g��m(�t�͌�+q�n�S�`����g҅Z�/+��ș�k[B3Mb��� 	ᓌ���+�DR~>��c�g�o�-�6N¥�+�M.t̞��@��ⱶ%�8��yy��_#��4W������V|@��g62��>� �c/ɾ'�ya6Nҹ`G��goT8�׫�qY���I�S�)6���N�m�W�
��1�V�4,�%ķ�w��L��T�(����љ��|?�/{\���~�>I8���@!��$�8i����X������V1��#n�ON)�I�y.��������ԙ;n�P��3+g!&��&w���Y�f��`����R�:����������E,�:�"�.�ZI
v[��%�~��o�1�?vaLD?���$O#�WH��$��[����Ze&M`z) �Oc�6b�D��@�jkt��g�6v�=�Z�L�wMߚ�+����cS'`ȳ�=�B���d���RFf`d7Zu���I�?�[�1�1��K��YX%�2ꢊ>��	���F�ln��I�p:.��`� �֊�g8���>BI_���ձ�8���!r�{�֡�d��to����T�ӥv�}[7yr��)�_��2��Ń��$����n��q�f��4ǈ�4�_X�K�x|�7hz>�F���,���/ֽ��_�	�hݿn8�#��Us���n�������ִ�?$����dl[5���8)���
ic�b~�)��Ȣ+Sn<�ϴ��~r��:h=����џ�s����y��:�R��ʈb#.��YAU�~�t���n7o$q>�W*&D�+W5�6��z��$��[`9���R)�9v�����*X-m�b;ñ�.k�����K��.�"�W���_�I�t}�?�zC��	��7: 1��K�6���S>UJF=-�,j�h�;�ǋZ��[�׀�����6M_�O����z]*��R���w�FJ\/�9���������u,H1�p��+h �Uv�넰�*�?�l�Y��-����0y'T9�>I�x���G١EUE�s�扤�����ɼ��򗫗��|�ܷU2���	��*0�W��+�K�a��U��I�f6"_hϓ�R�|*���ƇȰsZ��p�����E��Zs���ē^��|,U5��Y�T<��%
��u��]s�HY�$�e4ٵ�9����5|��q�O#��y5������ѥ��/��[�^��2k�R]2B8ܓ2���}�Ϟ�E�x��=U;�6���yKI�D�)��Dw ���QOR�����ژɨC��kt�
�zP�XK�9�襇w���r~sCgR�XQ�}C��u���`5e3k���I�|���K��H�8r��ND��v�\�~���a7!��sM�@��TX2��Bv�u���Yn[�続�jr�+��67��G�q�G�K����8g~� ��5��N,��p鉯��8�Ǻ�������U��;E5��۴*��<:{ 		��
Q�o6`�5i� ����b|?i)<�V��Bc'݀g+�� ���Wܧ��L�L�	�8�yld�$Q����� OA����+��-�Q��<�8�O����-�k� �{�R���i�+�5���T/�X՘oR�-
���R��x1bF�|��������埢c�;�x�a@&��8��FG�8Ђ��u���1�Xd�����\�ޏNF��ԁ@ۼ����7.}��]�$�*�o�bܔ8y.�"��-r{X��!�ÓE��C^�fܱZ��A������ݗV7IvF+�w���4�i�\-% ������%'��$��|��Oκ���%5<��� �u��P�`��kg��V�v1Y;�Z�~?D���"a>�9�#�o)9d�%�Q9�Nq��L�<˩2@2<Cj�� �<*��ϕp��DF���m�	
D����ה>�Q�w��8Ñ.��Q�;�玴M4��a�	�e	�`��\�T��]ag7�f��ܬy/��ʔ�}$�G�5�	c��о�Q	������>��9� \�5%�3,z渴��i���k��8`q�wĲ�t}���,�	}��a�y��E7�#�H��;��f�6�d�	��տֈiZ:�g(A���6dS?�ZRJ��V��l=�5	���3[7f`]JV��v���aj��7�����^� l��ldм��K���2�a�=|"[���d_(� u�y� �V���������3����9�%��^wP��[�Ӡ�i>���[����~}7%��#������|p(�W.�����帒�|6?j�We#X"]���T+(����1V�
\2�r�G�%�_Q�ީ����H���6%��%�lM�������t[)�c��K;���n4`��srB��������;u�:�Iխw��
�W��_n����k8P��{R3ޟ�h_��Z��ת-����pÞ�YR�ѵps���8E&�7�j�YǆRP�?���E��Č$���&���pn��h�`Ў�ƕ��9����dΧY��ŀQO���K#�&�D��iw�
ԋ�������,aU{�$"j!��4�r�K/�I+)]R��R3��/�l��彮pJUB�������U?�u���W�����h���&j)��mg����Q��ES�������{�1�6먍&���L�9zO�]����9Hu,o\w�e��/�_�1�7�s_����Ǭ�Z�l�K�~z~#%NBd��/{w�)��J�t���=�.b�5ô��!;��q���)���C�bߪ{g�����t_�=��-�n�&j�R�������@�Q���b{��O���%��������9%v۱N��j�{���]�6�բ��"�c�a{���Ò)��Y�OG��1����Ƙ�L���~�F��w�]"kX}_�mO���`ۓ�dj��)#���Ԩ�e
���C�#��ō������xb��1�T�@_&�׭���rQKF@���R���ezG�G�*{�_G_�,�U��o=�e|'�[���E�q��b%�]"�Ti�1�2�;�A8ghohjv�DPcv �H���+#+�F
�� �e\��@	�$�
,p|��#{0V�k�>�:�_dF^��R(�N��Cl��ݕ��a�x�}Ʌ�2���cS˺!O3��f�{�~#뵮&�'�
	 ��FH� vkB2�W���z-3�7�yk�w�q4�N4�w{V�	C݋'�w$�HFz�d����<�Ϝ��Yq��U|����Z@~5�[��^a��0�6�$�;�7���	�z/Rb���y�DKR)7)��哭/{���A�ћG|����v�dkr��Y��=����L\�B_�2���M�^�� �2Z��ӡ4|�ja��D�m�uk9�k1P�v� tUk�+sm��4U4غ��B�b=T�	�rQ��Hn�g�l;Uz�gE�d}]���P�e !��Jk��cZ�N*�r�]�Q	G-�`M��[;'��٦4z8���#�c�X}8b���r�V�ҋ�8A�?m��.����C�*A���Sy��%��|֌���d��*�y���޽��z#WR	��\xj=,$�+���BleQ	��v1�&�1)x����K7$`f�Cu1O���M���9��9�6IQ��g)x�f��,|7��D��_[K�}����zR%b(��z�t^������;2�t�/�g=������R�s9�e����Y?���m�FFZ����'7���{�U*�s}\�w�qE�y�'O��b�m<��V��ݗ���pX
�Ё#��b+~���c����6z���l��n��Ϝ/� ¯��[����/(�!U�7Vf��up<��2��g4-���'�{$n����=�yRͲLT#��NÂ�����$mh��6�f�D{ĉӆ��*�9[����h�}[�U�J�� /iKG��-K�R>(���`Ͷ����.g��{��btĔC5�	ϱ��U�Ĕ�[�3[>d{r�%��+5�PT����ao,y<@�_�T.�J�j-�<�g;������O�X��h��#B�?��>z����F�K}��f,�k��� �y:�+���>�GkѲ���$ؾ��M���f��Y�
,��Du���r��O��)�}��Nt�T[���0�jb@v]�*VϬE�->:68'�9]��⹜P�;�e��aM�[����e+��7�Ax������C�{&�)~+1�kճ�'8�,h�.�\�
�ɜg��^�D���Q�"խ�pn���9�w��|[��{�?�Z�Ku_DO{�d��q�!���J��y$�{�/eP�x��m��&\az������j�-7e��#�JًS�"&��Ȣ�yv��ӣ�~>���h	��y�z50��AR���Z C�Z�A�@��MI�8b��9&�D)<]�.�5olA�˶���e��6�km�4��qw��c��!��v4�Ku�(h��ap&�}��q|�^:=���(5q{��)��k����a[��g� %o:nX�@щ�q�y.��j&�.�z�i�d#nNf�7 '+�b�:�m��m����5��gr��z����Ϟuޣ@����j�^Ws���L�����b�X�(kT��P7�Ʒf�'�Wα��;B�ӝ�<Nu>�*@F��4b�G��d���=�x�.7M�8;�oΩ��6~��sHE6��b��Ʋ��ic]�dM�R�p	�m��`pa���N�Ȇ��J%a*�;�w���d�=U c`��SjlW�M��}DU�����rO�S�O�3B ݎ=K=�QV1��BJ��'��b"�5��&7ڤꬲ�a��Aw�(����␹r��v��R^�, �������7L���zF�↍��&�y3Я�� �����eZ�lu��(����n���I�ݸ���~���
F�o�A��~h��
��Rt_^oKw��GҘ�&J��m��d{���"��|�Q��(��
����`��Kf6F��mp�I��~)�Y_)6�<v�����͇7yF ;Q�~0$l�Hǳ�f���1�9��8�`_<��Ȱ��Z�-*��Mm�]u��S�_vq"Gu���!���EL_2�/�F��{��e��A���e��La�)��xp�Y��I㒘�:���W��.���X��i��a��i[�jr��������5��[��&M�r��&�F9
3�R�Vh��i�oI��&n]*�����U�GiEbM� �ݻG�����aӖ���U�
�[H�aɾ`���gb�V!��T�i:n߯��D��s}W�*c�E�g�o�]V"��t]��o�e4xʴ�eB͛/�]�PT��ru7o0\��ހ���(�WLf�x�_�A�(�}f*���\�`25�-����h\z�~Oư��o�?��� �!���F��|�(~1��ay�����Q޼���xA��ߏC��K�N2+6	k1���#xh�����|�Y��W^KQ�F
?�֫X%����� ��9I���b�#P�-]�������Y[��l�Xv�⩷2ɓ0~���(�y֞�?��6�߇w��̩`�VRl�I͛�"��eO�;��
��,��<p�܎:�FW�H�x��D.�����M�RY+����s����2@Zm�>�{Yk�A���K欧���j�EIv�bLI'���uY���j��}�� rx�6�K�G趮 3�6� (j^(���s%�U�����^$���m�	����K�g�}�µ����o��BzY�^��3�h9�Oe��E4J;nK�M����DT�$��y�䛛D�i�|�/�M�E��dM=��h.lN��A2p��%��}��\������W���q`���> ���a�XlxVHYEB    fa00    1d20Ocg���<֖����%�FCQ%��9��,�����✓��9���"	y��}��jp��>�20�d���l� ��"��c9l�U�X��(�@m����>���ҩ_A7��r�
s*E�u�ŖNn̞fkh��"�W0�a���-?��7��|�Ԯ�t���B���i���ںib��1��=������������.�<��b��ڑoc_$�Lr�2�h��y�p{ (��Nj!���|e�1�/������	�FG0��t��;�/Wۭ�Kܳ���m��I�s�7QE��V[]>-R"�}x}�ޜ/n��g0�L^H�BA�$U�-Jlp?��x?MS��?�洗��.����@�P���}WqF�HWc��h�z�,=��s$���AY�o;�T����f��Ɛ�×Ej��ˊ�s�L:�NE�+LԜu��sU��J͠��)Tʦ�1�vZ��)T���E
#��d�?���4�U1Ֆ�M��i�ѭڭ~��d7��c��:�P8�Ϩ[-��,�-�>��L�&�Kt^��V�t$[����O��d�I�I����w�mu��o-�MM�ʛS�ɫ��l�.���-<�l�k��J��eH��͒�8����.����k㒓��ım��YH�����#g��:Z:]�:��E��t�iC΃5l.bg����FP��W.�,�/�v�A]`��cA?�Qm�-R�&F�g���Z���U���f�ͫ${���_`�_��e���Eax�V���U\:������⾗&?v�x�;t�B���y؁wJ�&�	ק��ixN0Ұ���>e�^a�X�����J��]X煘������2pby%���R�v��tN"\��y�6� Q�1'(,�A�C� ��ַ�N�-��/���{������=]�?���ݔX/�(�Zx�c'��"p�h��ݰ������oH�J�h1U���Gk�~���Kw�9�ҳ�bɘ��HpU��z�!y'�|PO%�V"��!���Zi��h���X�9��A��%wDE����9��bY9%*�.�"�%Z%t�㝵n�{�*`;�~����"s,{���u~�'|�GXhZVN)+b��� ����Acug�$[n{�GQ`hp��ӌ��ţ�MX���@9��["�<f��ݲ#�%�F�,ⷄ��A��;~En�eLL~�]?��꬐o%�{M�~5w<�]D騾��;�,&1�QX]���F΁m����r<�/�����u�Ǹ��~� �Mj�	RJ�λL��thn%T���u�$��E�Uhj�@��^x������wc7�	���W1�\Y�Pޫ^��2���2-�q��jX�]��j8m�?���u�ʌ�F�}��'�mc��=���ӻ��F�P��"��R�r8�$e�8�;�S<
Xd�\���XgлZ$x������$]��^��m�w�u�і'����D���c_����_S?Q��)(֛x\Lc��Ế�F�4�"u;���fD�������#)�B0�?�_��0��k���~�qA�������$���-V�2{ְ�����g]8�dw���ߛf[�K�F���)X�g%�ˣYPZ��9���~k�PDc�Cx���ˑ���e���E.��A�uq!SҤ<�|�&D�P�۰�ӢX�c�D�WF�$�ELG�\Õ���	ë���*���Z� ��
^��s���ql��LO��q��h���x��ѻ��?���6�!��M��:g�9�DZ���$ys�h���J�3�3B��V��[��U��\���' L�� ��$�;�3֒нσ��
R��@�bL�Ȱ.���=��߾̷�t��؀S��ܗy�J�"�!��UO>�9/��b $z�Q��|}�K=����_
�g!Z[�v1���#�A���6��k)��sh�Ĉ���ކ-#���;�A�U5��{Z0�T�X}�{�_�/���>tG�|����j;<���-#������ ����oOIn��㔚j����,s�ݟ��'��h�?��и����r������[-�� 5�pQ���ݸ���1\6��1��ú�,�P\ݱ?�A���b=�Cj����ı?3?O��V��U��:��"��'M�ۤ�=ئR�_����~�Ԫ㲘���w{s�k臒�yC��Z�{�]!;���rB(i��[�m;���f����J�'�Imf����2K�7QԴ��ݏ�����;՛Y7PE#fĆjݽ���4P�,;��ŏj�w�����1��)��>4ϹZ�I[�Z'W^u�-!��͑O00��Ya� 捋�]�ƆWS��V�8��O�P�����\�a�3��r5�Ō�j�V�"Z_P��tA�@��&�;A�f\%>�c�������G��=G(�Y��n��n�@���y�g��2ƪ=�VO*�H����w�4_�q�ORpK|�3��E���wC�lB̴���>�0p.�p�bpn�h?��z!'f� ;�}�86���0����.X<W:���Ҫل�K��)��B]3���l;���aj[��s�{�,���sY�ki�+����2�5&��ׂE���V��.�7-̌4�:fյ�T0���R���݇�l�Cb a�oǯ޶ԉ�cS݈��g����c�4>-W����n.�2�wT!����[:4��8��9�/zVm�\�9��w��r��"��M��S����<*b��{�V����&�F�*|uk(|OBk�?j=����G=���Q����,0u��$���#;���i�܁���h��7�f̈����
}=�(�ŃzC%���D��L�� ��Ϡ~��h�����z",(;[ȵ�^�����Ĩ8�Zm�u�p-��S8�R�8m�f��e�^�t���w��O�mYs� �6�#��bmZ8��\h���������>�Y.���$-=&����i�},P��y f�炚�Bj��>u�5��A�k5��G����M��R_+�2�:cknG5Y)�x���l�8��}`���V�'����^�+ȩ*����4�j�u�|MIǨ)�;�@�_�P��Я��$q:ѱ!�ެ�l2��D�R:a��r�}����?�?��D>8� %�VKFo:s��j)��5��s컐� $�W��KMi>?��OR�R���bv#5��H��4�Q���uė1��D��j��=��$�̙Z$�la�U����k��ڳ�̹J���ߥ(Kǉ��F�ta���0�/��"4MJ����;bc*��nN 	� ں��q7���
�g�<��� ��
�W<�s��
����8�	��|0��!�H h���B�5��_�XW����������B�Ԅr^�H�+#��Qýg꧖6��c`j�X��g��n����=!��R��p���4����}Q}�,h�WA̛���6?>P�	�\����܇U�Hq�3#۾�By�A�*М��Ә��f���7��I�G�'$�WO�����5� �t?����%��.��4��V����D����hvw��`�$C��>�]Y��&���Ԍ�x�-m��^����+�]�p�br�*2H6��M*oDF�C�F�����';��Ԓ�p\xEI���R<���t$?1��ˢ�.��ً	� F�ifr��M��`�� �U�X����h�Հ��8�+��SW�+Ti<�#J�T"�j��g���W	�V��W|1���z�����1��kf��M�3mV��a=P����/hML"�^�ˍ�v���Z����~�j��p�#헟�!������%�{>9h+h��>ItTh�ˆ Xv
h���i��d�ڤ�ڴ16�m$�M'�;z<��)��6�Z9��@%W���jF��଀8<���"��NMw���.�H�$��`����u�j�E81����z	i ��m�Fj�*�g'�=1o�����3�_+/[���ڢ�"Z�~��0�$w9��K�_U#d�i�L>�97�$��+}�,+�~G,�,=M�F�	�,�K��M�ߓ�'����}���mU3I�M-S�Ń "����t��.�G#IKz-g�h+Ӗ;�KS��G]#��"?�vu�̔�k�t�d������K����^N�����&k����0�<b<��S�YS�WK12��"����8R�%�-�w,0��/�&��N��y�H?�5d��5�|W��A��vI@3L���C}�/��_ϒ�"��mt�?3.?�EdWMO�O�rO�j{��x�r�F�}�kc��������D���䔶F�>z4H��5�����B���!��\��
[K!�s��4x�>1V1�@�ƞ��I�$�
8o����[;�n�r��=�3q�z�R �Bק�C�{�^q��4n�{��<��_UBvG��G�)��)��<�����ŀ���V�O����|��e��fd'��*m���yʨ3�J�%[
�}%��ڞ}�d�D.���	F� N�c�v�yp A9'��V�g{���!]v�y2f��d%�?e VK1�#{�,	C������/�\1���/��a�0�F+h؅�G#S%gNX��\V}�����?�Log'�:e��Uu��r�f�~B{<�rQSM�����-Uϡn;�N+���	y���}�4���3׫�-��7Fs�]�&�1<���U�P�3
�U�k�<0�՝q70�DtT���M ��EVH��Ǧp_�M�ͺ�>u�?`��]��U�81a��Ui�d:_p@��Ô�GtV��b	��C:�d��:N��B�<�	4��G#�G��,疳����z��	sR���3�ى\b�}���-hl����<��iDO$��r �M�����=F��0	0k��=�T9K5F���c��|r����+��~A�&xQ5G��2�m%aU�Y
3&d�\����g%�B�P��>K���}k7ez�'���*�Ԙ�I<%���0yQN�fgql�dPQF{ �G}�����:�2c㠭B;ËX0���VZ!K�$��\б:=b��[�׾3D�"�Ġ�����i�ې��-����l��\eJ�NF"��T?T;VJ�% �<�f�>�Hy%@.���!z[����I�����6�}���,0�e��$�?�ޭ�ٽ�;Q��9-�
�MOid�)���x@Y,SA˹Į��ym}ʯ�A�����L�p��Pl�f>�s��	�;�t
{N��	8h&bʿG�܌T���$�>˳�������~`ncj��m��4�Sx�`�6�,^�]���7J��j��5	+�����m�}��� �	q�����<{EQ9 @��*qY�S�b�k��Uk�P���N��s��T�ͅF���330�Y����]�<�LVu�?F�J����������c+{]��ө�6��]�=�����D.��=����u�Y3�Urm�eͷ)�s����)���G8��5��J�τ>qا���\��?���+��=P�y�q<�WI�K%�Lԏ�'����!�Q�:q9*?ɉ�EH~�i���z�6V�k�,�Z��«���%��W�3�m�CP��o_hγ3����W7���m)JS'\�KbUճ�HY�z�opRo�E�3�Ԇ?�(H���R�	a�G�i6��z�c㜭�>��<�|`��ÌA~���01���&����֧��?���hB/5L��e?�6��0�J�u�|�����Œ9&�zMBA���6O�%�421�ܕŪxK<]������V���!�(-GZ�|�.t�6��y$ED��6���Z����XT�2�E���䮅��t����An8��Ak�4>2٥(�F�abB���C�{k4�ǘ�%�u��P��VC�|:Oyoh)�\ d���U�s��L܂9
΃�u]˿��'4d&���e�����$gP���8�4,9|q�(�t�'���,���2��wto-�{��'t��S��4��cF������i���W+g1d@��V�j@*Jރ/��R{ �\en�Ȫ
k��Sg��2e���D�9��I�l�^�H����O�Uo+Wm_%I��cRa	A|H�p�Ź[&�a@��%ˇ�W_gl���v��ޚ���z(k�C�eNT����6���$ae�pV%t�S9��7\��!��}]E��]	t���i�S>U�z�T��`�%)� @'(�A�A�1�<�l�h�4j����o�Ӵ�̰��L��	�z0����[�Wy��ҟ������+[��ȤN���e���`*]��9��"�#�G��;!s<�++��i���VkF�����6��2�2��@D��W��kk�T�ܼ^�&�v .��I��$��P���u��n�o���-݋��ts���*؝��) |�Uc����qQ%��D������S۲��:ߜO�*\
�K��k˘���EVb٪�&�b���Sc�+\�c�L��^�Ғ�)/g�YȎFľ����Y�vq����8S� /b?s�'�x���$�Y�)9�X��;V�M�yp����|o���x�b���D��ߎ�˿�gB֣td�
OM��MM�5ȓ�Ak��zv���9�I�����W1x�ڇ� ����ߍ���]�X|&Η��+;�]1@/ZvlxR�o�ɤ��%=
枓5=nT�{;��5��;�C�N�1���.�1�7_G��n`���]g)R	'K,��F҇�����)l�.&�\y��X��U\�Mgo}��P�&&P;�i5$��RݝfA��k�������L�bǾln�7z������ح�����	?�߫0�N����j�x��V�N�a�Ğ��:<�+~w04ϟ��?������*3s��7!8��|Wb����(ʠ�����ǋ��/#�v�b�2��x~��2ג�x�'I�9ͱ��sSCJ$.^޵��4�����gA��O�S	|3����`�7�w�
Iiw>:v����E�у& Mġ,��C�)e"�4̌�����;���'z�9.>�z~9<���<�D������fh��"��ߕ�p�Z�\��������0q��w�v�����~e}slk^'C�콐�L#<1����e��I�8m<�T_~"�y�j��y<]��Zu������>%�|�B�P]T��dF�x��%�.X:�7��J.� �+�&����5qZ_���	~+��h�B��
s���I�N����郘{�p�]F��*[���H��ڕ�#J�}��A�P��%����p����1�= @���y�(�tҵ.Sx�{A�E���[|k>�{�����i9�
�ݘƍ�,s��8�&SE]��4}C^��OO���P�h¿~Buu�%�G_��_T����SC�xN�x1�\�	o�%�XlxVHYEB    fa00    1dd04�RJ�����C��ϥ�H�E�Tp���%��um����1^9F���$����d;2��E#���CY-;�wb>G�D��a�_�_�-f�p�K��N��� ��6�}�3� �F�QF��.�+�`R��X��	�{3��aa�w�Y��}�: ~�����nXĳM=�K�����f��E�H#�e����Y��ٗ���j!u��T��4���v����K��)�-�s��Y������cM1e��e���v��#'uV�@OcT���9C 4s���~�
�5�t�/��|"͐$y�^��tF���Q����s&q/�o"�t�=CM�!#Nc��9��Z��%AǄ��+tm����+�����+않�t9��̴��N�hW$i�
���WX�)�0e������,` ���`�_�������p��(.�g���9Pq�i���X�U��{�	�H+��8�S�.�ئ!������ޕ/�l�0X�R�	���l�GMJ�%$W�0(���U^X�{��W�0EK�3yf.4����*��S�=̛+G*��P�&�zJ����n���%��ǳ;�:�U_pJ���U��4y�R~�FHm������2͕<�ܬ�9Dl���/����8�U�H&\-C=w�i]��I�B]���'�������H���s� أ9Χ�%R�!=#�:VJ�t����-P�k��/��E]��Q��bғSS��w����	imY�%Bb�5�w.���'�z�K7�=��,8�h��M���T�]�`!x*�c&������1{I+P[k�z������,-��j�`��/������Z�c®�9^\� Z�W�5�
��m�����k�a����@��U��AU��VL�
> �Ŝ΍D3��F|�K�^C�H���28�O榢���M��Z������%�5i��`w�'�I���E�{=�m������*)������x��D��=8ȷ���E�7i9�1�MM��c�Vs:g���ֳ�5�R)�緮��GK�i(y�4.h_��f�k�gh���	�,����ksMF;i1>��T�ń��	��8�R�09Pµ���!�J20�����'�4�Gò�~�8C�=�����\/ɐ�;�8V���$��� r ���0rE�_�̘@��|<U=�(����B�v�����(x�wl�=p���oZ'ZQ�����Aq#<��o��"�1�a�[��G�f=���C(r�>­=���Bl��,��|��iyL���(�a����;t���i$�O�vA��-x��W�̻�T���e��g�{��w�!�Xy��bUɪy�YwnA�#��ٲd�(�
�l�D:[������������B���EC
��?^�Eg��i�8�����D`���d6{x&��lI0ס�*�X)bd<'_~RO��4����B���(�#ZI;;��0�9id~���a9�f�4|��s��;�{�j�"���r���A�UI�����0�,����1S�r�?�6=���o��!� ����|��Lg��Ǯ}����nS�F�Kω<��Bq�5ޕz�KP �xbI۸���&���i�緢�8Xwd�=A1�*�ϟ��BYʰH�Ù��$��a�#*(�2�;�2�QR��wgc�v�;�L�?��chk� �Y�cD��H�����ks�2Es'�#꒾�!��ri8����[��j8Il�Q:�M
L�Q�0ߗ���|�*� �OX�f�s"Fᙯ����7����+ 4_~e�}^E`���ݕ�g�(1�w X&�����!����+A��^a~t���6F�h�{nE'/���~�;�e���ʀ*��,�V:������և|,`I�\{���k5���������g�@m��$���Y�{b���Hw?[/|VE�*��xk3qUA�Ӏ�(
w�����E�ZKAP���I�l�-.҃ �cPZ����oDK�S����X��9�s J���II����S��uU���ҁ�պ��e�u���q����ʜ�������͵�b�ì�º�+���8a|k�iU�d@���u�x�0y�*'Y:S��.�N��	L�_��y���'wa�
#B���+�Z18�H[��b	��)�T��Sɗ�4>TjE%�HxH$ů�g�h�NVE��/�80�Ƭ0U^�P�0�Խ���y�N
���a7�!���wp���;eӭ����Y��|�P�0�����$p�{������P��N�+k�{D�i�����ug/B5m򺼟�lw$U�\(.��6��CHM(uy������P��q��Zir%�ZN8����&$JP��M�g��x�b� M6.�����ey��~_h~z�K\�c����}P����3[��D<�T��Xi^l�᧢_����^k&y��y�y�~�R5�(�����ǉ)[��r�"��.��7_�n�;���������O�l���xA�:ӎ�v�>�D1(�,�V�	'o�1"�O.9q*.d�����0H]��5�m��?����5X�z�Am�һ�D	��5h)�z�ZoGS´8_~��+�o 9��}
�Ҹ��J[23��׋�������%sC&��@J��G�4 ��Ǣ�oZ�������+ה:��w5�҈���l�{�q������%JM[фM%�nƻ(;��2�Z�����R��LB������\b=��:���JA�_^z��Ӟ�$pt9�F��o�ފ*����2)�z��ڣ<���CK��nE�_�Jx"r�ߒ2�z	w4STL�O��B?�dJ���t+����6rS�+L���b=�ȿC��>�����4�h�0�{�Qy�������OV\O���a��M�ʥ>�q['�]b�����4��4�*г���)c	-D��/�	V�'�1��*FLI�Σ����E$��#@��S��ā���B!]\�,����J�&`|1u�+�.ݍdxNQ�w ���^䆬��GC��d^-O2b�x8�:��(�	�{��@�Wݾ���E`7k^���DÖ́��Rɓ6U���P3xNr��Y��R�5�9���=PX9r��� �>��1�U-����F��a�"���p��:��~��ݥ�EHǫ�Рff���V>溜$	�:�g�D�I.�p�!��_�������}y�&"�o:�#`�2�7�i�@
E^�6�U}�iH���~w�5����[��sa������:�W�}�>CN�/�\��y�᭿�>:�Ռ}�s*���W�-9Swa��x�\�ԭ`m)n�^;�z�kP����DU�kn?�OYX����G��~���V�������O��2�)��S*�QD�h �����$TS﨣�H)@ЅjM�5՗2O-!t�妧�<�c�}��F�=��s{&����|�ꍅ����o0y������$n5Zs�:32��m���	'oG}j.�92�|~�#���%�'b������_0wW\�v�_�$1y2�ѫ*p¸NVeUQ��*_!�Q��ú0�֐��_]m�/nm�F5���S����<��p}��������8J�w��}�A�7�x��������t���e���cgC)���+��e�+�n&0*;PX~�ὑC�iT1�ḜX���S4��V� �P�g�?�|Np�NS�8`n���7��'�Ȅ~!"��L�x�����2�U!�X���k���'56ɝ��:�~s�n��	[�G��F��6�B�~p����D��pݟ��Č�D��iXa�g�& �d�>� E���9.f�-B5;<�������/�7S-2�\p}S������Z<uQ@y�Zt�ezM)���;�^ �6���=x�ҽ?z{q�뛄��V�mU8�)_{�+�<�>�LU�0|�f�{e=�����OY���>�ƿ)Ya
�vV�5�[Ͷ񭪚�~�i��O�����nz.�����Q�k�N_-MB���;)`ܐ��Zq���G�k�1�t����|����{F`{BJ���4��)�b�-DgE����w�����_������f0
`��@v�/R�S`!��c�p��8�۪���	P�K��9���*�*�Wjbb$h���Oa�5#�SZ�z�ǘ�p(�Y��){tX����ݔ�
�<D%f-x��|����S?U��@0�jxB|ܧ|�N1�f]���<����B���ԟ���
v��61������c�@�tY�E������C'B��Rπ�q�C�8�CUˈ�7�`��
�i��ؽ�r��T�����h$���(�
>�!�xR)���(�)k�K���J�Vl��3&�;�S�6�mߋX�~M��/��y����I)D�X~���®R��+Of�.+e��b��.7-e"�{,�h�jX�%e���R���CY��Y�z`�[RJ0����V�$�|!��X�-�R]N�W�d��t:�x������VO\گ�]���Q�~Ex�8�%^�Γ��k�(:3L:hvdC�B��,��/f��d��s-���<���.x�M,4
~��T|z-�R����;_ ͚Hm�.��Hq�����y�%�.���B5�yS����]����Vnj\���Q/9�˕vc��&�IE���꒏)o�S��s:��d��<���	�_�]ל���),t�h��o\���A���V9d�I��7��x��̂3%()�Pu�&A������wgsh�p�B!��B�[��8��}(y�F�)r䁧��$����ʁ�L��HzU��s�Q���ZN�S��p ��6�ZW�ƚ���4�@@�M������?�����3��d��̼q��e�g!uȴ�xݒG��Ƴ��k۷%�Q
���9�����4���N
�BѡKjq�Մ�3'>:�^���nd'���<n�/c�*0$�H4��E�ojM�/�Bf�E�׈xa���0#��S&<�ڑu��j�O=��B^qi������	�P�4c/,�)�u��j��r�L�$^/=�|����M;>��?8a���M+Z(ʜ�<*����XJ�����gI�q��n�0֭l��[!��"%����A�����Cp/
�	�i�랔�c�t�K������Sl+�ԧ�K�m��G�Z�w�i]�k\�[Գ��ݳ��w1A�!Q�k. �x�IW�5���xc��~$�u�$�r�$�^m�xLBQ1��h����*��b�Q���E�ćzu0srq��u��������ڍ�����	Tڽ%���;�t�G ���j���<�΅��K��Q0��B+CA'���	+4;�U8;C�w���BCDD㡖TZ�����4zP�v� �&�ICSK�7Ē�Яm�#�X2�	���3x^Ϊ�޿j=���"�\ݧd 5%���;y6lS|j��Y�&A?A$��&q��\kG:-j�a��Κ<w�p�ч�6(�h��p6��L���O�'�Q�[�IWzWuZ�@��AkjP'׽"����?3��ؕ�$�px�M���\x|1+�;Oqm�79�2� {�Xh��\x��_�{ڎ�Z���es�߸�7�O��L�f�<���Ӂ$��Re�[���#Q	�y=RR���#��G�m�,�c>_������G��ȕ���S�4����|�E�S���x
Q��K���E8���u4��&�j�qM�*��i}uj`�d;A�{[��}�ͬƺ7\^]>j&�1��MEO�0�~E��(&���++�p�Y��E}�>�U�+�.�|� I���vݶ"R����T���0@ �V'N���>�X+��R��bv�K�zˋ�8tޓ��p�����؇r:^�kB�O�;�c�Q�oõq�}=Q��N��Bn0~N<G?���"8F��BlJQ�*�+:�Zd�[�2$aMKF�ov���z��&��n�Ý��,g�.�xv	�.Uϣ��s�\���n~j���(vAP2�E��Z��\�¸S������G�(��{9-?u(&s��w�jb���+zXO�*� �>�#}Km�;�Cy�u� g�m
�R+�t�`ؙ��u<\ҡ1GD�>�\c�pX�{!���!T���=[�p(��b�)h���ѳ��5M�5wP�?�h�Q�1�;�Xc]�vuET��)O�|U{[>�X�)4�L�I�Eg��R!$��q�/BH[�$|(��sM���x���UI�|p_��m^� ˅�)P�c��[����Y%�Lh�A��o�E
i��^����\�fG��*�L�,M���*O7I�;��v�~"�"^O�'1u��6�A	sx�d8R����|OR�����A�����4=}���P��5ɉ���mTY��@e��4#��� �rA��� �L�Ԁ]˯�a�'G��3�s{V�^�i�`�z�l��yu���k.�4.T�����&i�O��x,ڱt�\[��^�Α�s}~��je���|��Y�O,7Τ6<x+Һ����t�-���j`*�C4䨣U����V1���2X���!W���Y@'ie�,d�W��$��-�m�n�Mf� �{�ul�f+�Z%����tD��a�1c�ι	M	�VmP3ۄp�αQ�sS�ا8��>?]M�_]�x��YݝD���"�Aj"�]R�	;K�|�nUZ��P��=/X��B1 �ڞ=9�y0$���&�?�D�ջ��B� P��Cŕ$ ���m}���P�oy�}Q��N���<L��;	r�;�QE88��b����t�f·{9� 9<u�/�^��\�l��(J>�zV�w���޶���'���!�R�	ԶoR�LC>�����{o�����m �������vH��@�c�3���5��j'�#lzG"���_��nS��HḰ��2��u(>9Wӝ�5y�&�3l��jDb"x�G'`�t�nP��嵅ܖƽ@�N(�)>yh�~�f��WsɩX����1vg�;�NG�`�Y��Gs+�fS_b:1{��a�Ɖ���̡Ej+&|�("Q��s��;#2v�!`��/�ׁ]�T����5秃�B��UZ��X�X>���VZ�N���q�Z P`����g�v>?_�z����q�LK���B�4o ��I*]��^�)O��V�Lb�vQ���
�v�� �\���׳��F�T��ߘ�[�-�E��ڢ��`�B�
p�n�d����PS�T�b �/UJ.a���p)����p/�h�K1)�vr+�/[_�	�ox}U�����xCϘ���u�����zm��z���Y���w|V1Ά{+�\Ig�$;Lv�];�2c_uW��9a��m�@3��ao,$�[1oSp�	D2ۏڗ��ُ�����K�j�)�W�W�m <ԓť�9���.[I���rs��d��[����	�/P��;��\�T)�%��~�ޑu�wy.,��7�^�^�ʦ?��xC\���0�[^uc�XlxVHYEB    cc25    17c0O�K!7�H�ye�i|�g���G��N�V��쌿�2!&���nBdR�|��T�ë(r�d˰����s�W�kZ�����Wm�m.�`$���kܙDm�Ĵ� �-3
�^25��hmO���l̇l9@Gx!���/�"AIm��I��Y�>�ƀ6�;e;��ߓx�6�B������t~��ɚQ�l��5P�j<��2o��tx!wB�}�e���Xuy���W��Ds�2���}�B��Q����j��ߍ�)즕-0�5�?5�Da����X���7��YG�+��x�f��/�7��Zm�h��%�l��Z���h��@�z$�a��hN��d@2�,&���'(�gO.�0���ɺȯ�jUB�{�����~�Y�-z@&n����l:S��\Ê��?�9(�����Rf��c��c��kl5tٱ'�`za vL�X �O�őV "�/?��U.�i�@at����Z��ʄO�Vn/�-k������x����<M,X|���@�C�\� E�8���Hѝ�}5���atHwx.�v�}q�`'D<J������l�w��*F V@\��ĥGv���DV�`�L��QN ���7�-qǊ��
,z�Q�_�r����}=�j:�����sE~��ޤ�I�u�Df&
����RkcΌ�
9�nTY��"���L{�������B�m2G]�`"��#�!y����a��/���[:��i�l���e�9���w���k��!���l<c��q%�C��T�h����;(�q7^p{�H���۶��ԄX7�OS_$�B��\$N	����,�a�W�z'��O	ֆ@���O��|��n�$wuw$��D���T�(K�;QL����*�5�� �N�8YcB�bMQ���д���e^�I���Mҩ��Qi{,��n!�͓^�E�wyZ�Ç���R/�yCQ�݊��Zb;5��,ɧ��#�A�[�=�m\ 9 7w���H5���S��]�$��>M�����5�W���	����җΐ�Ǳ�w�u�=,�z��נ�����6�K|���\�����!���@�l��H�!l�͐�X�rM_��w�|��#�~�kn�*��*�fq��K���q�9�O`1h,����2L��h<�i�9#{�R��wھ�S�%]�B w>�3jܹ�^f|*��r8@w{�=�^��"�V�[����Y���q��;�u�ksG-c+i�$Ke�D=�K����kl�6jJ!���st��۷�FO!PH�&�0��g<p "�S9�{�75���R5�c�:��*�*��!J��Uv��n_,�E>��3Nt��M�-��)�fz�ʻu�x�4Xn�h�����v�UUD=���z�Q�@Z����I!��h�m��(p��o���>E"�*�����>�\���� W����y�4�T�4��~ؚذ94B㝑PI7:3.2��b.o�U#7�����Tw ߁�����JY|�n����<�˸����	�aPi\6�����������Or�f�f,�^O<r��B�Х���1mwkh#5�<LbDl͍$�!��b��*Gف�c��]p�|���.��v&P��Z���Y�,�R~	M�Y:Vn�[U.i��=>Tx��*�!�Yr�?^��!��i�"Q��t,e�'݅�Zx?�Eß%;��8�21�xi[	g��h�uմ<�e6e��U�RfkN����֑4ɱ��x�������k�0�v�M�/��&�E�:������|���<�w��w�I��&�F2�u��� ���L���a@N����T��)���3�٩�&�d4S����mdr'��.]��g!z�`���tX��$$�+n� J(`�_8IH�I�������Ɨ�� �eKA/&p;�n�r��ܺ�:���Ӌ��@���ct�)���<~�*g�	f��|h�Gh8�N���]�ٶʅ�՜�жZ�!}��6��'� ���*��{�|ҟ��]�	�ƈyo��˞���PM�A����<�!�Qs{Pq���������u�2YX�a�&�f2_���;x�q|w���3.���w|C՟e;�ύ�t�N�D��,���^V�������_���+m<��Ӑe�q���͟��$O#�>'��"��2/Ԛ9�L��e��蕩_0ꉦ��_���H�H8���Y�v�^��ݛ�D�abv��f��)�&M>���@��%����Η8�yqGvPPҸDB���l[:��h�(.�2�x~Ѯ\n�׭�D=ۭ�؆.�xցJV���{����4/D�򨖚ςW���ȬY>2@�x�����anv�I�����=\AJ����-8"���3�{s觮j�l�_�Иk�ا�=�/X�pCe�j��X�y�z�Z��*c�O��ܖw>�I�Z�xl��O.�
����2��S�I浆潘L<c�)�	�K"��$Z�l]�Y#:�:'l��a���<��~��0R~���;�2v9p�@nJ���5����0Vص�R�6�HH�SF��h��"�/�\��e"�Ś;���=�
�c�$����u�Z�7NL�P.�HE���T(q;�as��Ƅ3��#V����w��k�����Q���9N�uY���3�r`ăz�P*b#XKft���C�Y��wɧ��z��1�T��_ކu?w�a>�&���e�i�N���~�$��r�;�eX?�����B@nPg��"��b�e��r6�'��4��@�i�l����0��~������+�)~�|Wú��n�$���v�%�e�9�Z02߷.3�1��kH�i��q�g��a�d_�O�X�i���/�<a�W�q���T$����&�� sҍ��Q�0yǍn��^��N��6��U�y�pe���i�� ��N���TMM��j�-��`
�$&dz�KWC�$���%X�N^�^�`c4��33�RG��� �@�7(���oڼ
��[t�뽖�j�mC�+fn=<��_�f���Si6`M����&��o�/>��f�g���M�o0�I�Aā�5��u��;����M>�w�S��yUB�GJ!�6�h2�N��":����")Z�.t�7[+�K�Z�b�����9Ů:��P�VR!��N�O�ټ��^۫w���-A�'Q�-U
�(Ň4���\45?;Am��x�Dʣ��`AL��~�, ���+�5[���{�Hz������I��='��M��T�/����|��g�FAGu[ы!��ʤ/͹d�N����ғA��QG�Z#|gT!���֦��{/Z��%�͆`��O���|�&�Ԯ��p��b�w̟�т�G��z�:���>������ޞ%�*f�`!�/ӳ���н�]��T�S@%R���$u����6�U��a��"��D.��bݒ�����+,}�\����Ǒ�?f<K�,���8и������';�f�/��w�|u���2G�1�nD/�a����X������:sg7<�ϛɵ�z�68g�Ԫy�(���"?r��#^����R�%���Gc79����H��Ƨ�P��[_�y�្UAE�!�f8��=t'����v�6.h��#��d
�`���?F�@�<TM^�:w�-&��'��(6`��,��*�D�9$���ќ3��axd�>�ԃ>��j�9���|���ػA�S�k�3Y5�օs	�t©�1�7��h��Jc����휌�dh�Hj�[�~[iUs�أ+�6Cy��o�χ]*~��9K�2�!�\����J��O���^�R�gL��BݖB���A
�"Y�<�-	�l���rE�u;{���G��%1nD=�����b��V�N
3�J���h;���?u/ͤ�Z&8%�dq����s�>�B��J�i�q�
���c�5|����$��[;��ߊ�X��+��W�b��'5$���>�#�^:�={���e0�d����j6�v1��`X�M$�.��_P<�X�q�݄�B�(�ʊd�쓚��;����������;�j���O��r�r4#7,�%ō��]}�?�c��T�'7x!���Ĳ�����P�g0���hb�)��kLiK�e��tj �ڷ��:2�n�4|��Ѡb
��@5�7�9>0�{)N�`k�0���*��^�]���&�~�y-�?L�^������ܫ�u�\�(a��{�p�T��yfC��b1�o���*�T�#�)�e�f�(vb�D�4u*E3p��Bv��bX�!�{Ø7�EZ)�N9	R��2+�)�5��b���'�<�g�N�\=ی o�U5���Q�u���������*�-U��Xpm\*z��70n W�ޡ��&�a�>���zj�ꤽ x%z����5ʁ�Fi���[��0/b��U+��5�;�թ&oD�8�=E%We���vD\��ݰ�1���Q�0�b�[���mo�%;88p?$�G�� �P
>�_�j[<��*~M��z_w�޸�������|c>FB1�I�F1��^o��w�1i�\Q��h9T7y� ��#'=+�й�nx�#�J�� +�O*$`\��z��h�~xL��m��z�$�#�iv#a{s�ϓ�*��8�FY�w�ja����\�[8W5*d�霜�]rD���0��a�ـ����_��)���s������7Z+�1 ��x�<I�H@����$F_��f��iv[P��[�װv�4`�^ʜ��_���l/گiR�n�=�,;s�1����rr�㖬Ph��w�i���)F�_��d�]"�\��h@��Y#�����]y�>
P�}�j|�D�Y0c�$��ݝ��\qsp$̖���<��g�MŬ�63껑�X��I�O�d_�#��q�6jsϕ��`)&��'ks��d%�Ğ1��(9x�ͧq@��+�8�5��HX��4Ϛ�j(�~u�t��y�&ʗ0�4R�7�S���j$�x`��c�٠�
��=�!̐��M��J�X���^��Z���#�$Cs���V���m:�I&��Q.@}qaW�Ҳ�/"�h�
���21N�p�E���ߵ$���{w}��8�fW4�_�t>K���N�yz��s���z&s�6��R��rF���6S��(��3,w������S䆅��B#��3�K��%�S뺄kj:E�iE�vN�r��̊)�p$wH_(	��72��X����I�^B'�XTQ]bJt�̄��S6�!6m1��D��s�u�.A@���ua���	�$U0�eIմ!�ń�"��b�ӿ��ī:��i�ba�i���F���Iq���p��bۗO�p�x������Yn���%��L�v�J\��/��8��`�`��S��<pۄ��B���k����?�z�oF(�T�uz������G��AG
����溜�� /�m��t����f��#��BfxE������]��@�4[�ɏzzm���<#�#�J��ǰ�BΜ �c꿛i��c[��tσ��6Ztf��L�2c�»�zS_�,י*���X��͊�B��,�Tû��;E��#%,?�%��W1?5�9��������_T,��P��/���k�Yv�3i��K3{b��}��|s��)`��y�J�LXi��
���)�we�K��r]��x�5g����ԇ4�t�_�ИܤQ�*��0/�M��w�����G	�3s��5�6��7��1�<Q��qy���V�yp�7x�x��r:U�����¹�$�Wg�����m+��:�\q���9	���D�o�i���5�nt �`�`��f�{���H�'HHû.N�ٞ� A��*��y;/b�y6���W�)�䵗�u��9���-X��$x ��W|�dBGp��.��ˍ�5Q=LW�_ȩ���]^	�>��vE9�,)u�����.r�$JkR+^5�<8Xu�F}V7��:���T�Ҝ�hug�uڞ�Ъp�˗�[fn������