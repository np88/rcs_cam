XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��)��/�cY8Z�S;���M�X@/�$�u�rڮ���U�Ԃ4��g ����d�?��Nd<��5ܓ�M�]er-^`�V Տ�dA�0��P'ʦ{�"�*��=��d�}$���L�֣Ӻ,�+�x�}�	�V̤���b�z�.c�h
HW�kZ��J����Qڵ�wq���q�;��X��B��b�&Rq�o.�4�"����vn����M=�ū�?P�s>���b f���َNTԸ��#�]�P=�{�Y4�-V�e����@vo������E��4�&3��i	�2�m����N��.a�І��e|t��VnKgU>�ѴFhœ�;��J��L�1�2o�t�4ėu�I�lBq�D�%�d�\��gĠ�z
D���8���b,���٬�h2���7�XI�(�>�!"{0�i	�d�����=����%֒D��[��u��R 1���+�(�9�MA-�U�j��8�u<,��dn��V�씙n���y�9Vn�|G{:����m|�	  W���M���~�����A>�w�S������&��5-�S)=-U1a�6"�;$t�Y+�Y�l�F�Ձ޵A���Ƈ���сk��#`8�D����6S\�r���d��r�b�e��^وu�@/p��y%�5���C	��Y�@����$$lF�<%P��'��8E� �&�
�!ro������5��*�X���Is�aׄ�	����������Fv��չ��i��l��d��L�:�zJ8� ���XlxVHYEB    15c9     860T�ij[bSnI+�4�����C0���V��e��yHװ�F&�P�c�N�o�ש1��D��2-%"�M�Qꚢ��|�QF���i�l:�h�-�u�3� ���>K����~�yQ�e�Ȁ'#i�-+$��� xZ���g��c�8�b�ܠ�k��$�"�ˡ$dV	c�����Q�"��C���6�t	E/�h�\"U��7 a�ow�O|8|zM�9D��?ഉ3Y���[��c�]`4gM�yL^9�j�U�]2m =��iϒG�
ef��j��04��|P3�c��uF�&��Dy��Bz�η
6;oy��鿒Z��0�K��)c�>���qC��b�w��`^*."5k�����������_F�M����+NDU`w�n3���o�,�K||��PPX�s�9�}fb�VB�E�5�R�aK�Y�Nk}U�]�q�r�ʺ�U��*~i1�?�S�tS�?6�P7ɟ|��1?h궼O��`mh��%
z);�BF�uB2/�M��+0o�bګ��K%�oe�L���]�����T��`���>e�ԕ��.��k;TTZ��
�͙T�}lӕ�w����@>�C��^١@�k""G������5|�Q��q��׶��֜�����m�;�h�M�fc��t�D���,#w.}ӕ��Q��c������A$����S�m
B��xQ����"�U���{R@�n��!e$U��zb	d�jt�.�S�ՠ�夽Y>�j�����0D�0D�\�q���Y��(S	���J���"��8�WG��z{
�R��GH4�s�Cх�`�"�A-5��Ͱ�`W�1N���_qt����*�VH�w��kOxdv�G����r���Ύy:'���C�8�>�@��؍,�/��3I�Ddg��W�+���N�^�j&#߾�5Xٓ#�[U�J*�3�J������rTW�`f����̣̤��ڵ��N8Y�#M9೑���[c��E� ���?��Q,G)')��6�Y��ofX ��Ssэ|Y��@Y�Łd�G.|�L&WA�׋161��H��11���v97du�>O�	8C,��� 5�=����;�1��H���\�����x�/�0d�N�n��Q��=N�c�o�p7}O����D3��?��i�fXɅ�g��q��w�(�����
«��}}`�6���_3�'�KXKG䗗��{�L1�Vp n�	>��}�6b
2�Ӱ�QL~F�=h��K��U�b��4_�+..EPw{���)��C�^]���>��e�_��������%��|��xC ��xL$���5tg�3z��"�.vj��Hvdw��a�!O`S �g8l����6όZ����r#���{7[�#DK:YG{�纎2o�{e�rUz��y�������])-�M"b�9�E���P��>(���V�4�4o��*���7�փm�I`',z-RW�}?�䋘m����>���U��:�`�;%�(r��\^� *uZ!�5�w��Pxyn�ݮ��L���Τ�T<�y|ˬ�A�K���Ba�]X��g�֋oYʤR�d�&Tq�:��!t����k�w`8���J�F�;���h�%�5�δ��Hű���:�q��"��{�!���^RtA�j х(B;����ԣ4���_)KW䧡�Q^�9�P�q�DtU���}����t���7>���.�Մ4�B�=Ia1.3�TN~S��T�KxG��n8�|[F�ɇ����6�ũ���f,���m9�X�o���l=�?����6�+N)v\^{�`��!�|���mO���*��4TѤ��8i�O�>�9��Z���Ɉt��i��D9K��QV"��xx��榈����0,����e���xm𣯡]p�y��0�(�%�Z��K��m;�tn�x���@�_n(�d����x�o��P恿�@$�e��O/�V�ċ8��)8��c�y�
����~��#t"N��0�`[�`�c�2��<ԕo����(HwR���[ַY�o���?'�����zi=����&��b;$���3^�ߥ��ߛ�?0'�?�=�1g�c֯QoDG�gt!�[��̅ pW-