XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���::�}i��<}'�H�f!��\���gIl:��+���ޝk��r�GvCSp?B���O)�Į�a͌�kD*�ih�#�N��@Ļ�Pd��i��.~o���R�'�(Y�<�Y��i7f�������^��Ypɹ���!P�xf����Sb+Y&��� �z�GF�"�Ѯ�"��Z9Ņ���8���G���p �Hl,��Rqhq\�c�}M[��e@=5���m*�UeV�����W�E��j�BÒ< ưԄ~�vz���K��EN<�����0�E*Y�0�m�$�2���!����Ӷy�X�Cイ�z�u2W.>Āb��+ʒ4W�s�+2,48����M:�琭����м��

[�
���Bt� %��l�օ�����s������������O�}.	!,.W��N1"ݩXT �d�&��~���}�O��4�8�᠎Z���Nd��s�.���o1��h�|�sZ�LФ��J����u��Ҋ��Mi$ ��<�Z���,�)^Ҿ���_�����hʀd��Bf���	<��؞�F����"ģ�a@�NT��HT~z?�YIy`\H�d�G7D��n(e�E��a@Ґb���Xh喔a�Dm�����'�Oq����ݗ����ӽi�k\�pc�_$¸��� ��<�-�:�����.l��
�q���q){��2��>���v����SS�b�f��&���ݱțjP?�!W�0g=mu����NXlxVHYEB    d7c8    22e0�w+� �o�Qj��J��Ϸ��f3垡�	9ZG�&{��Q�H{�=�Tx��/�j>ߠe��٫��|�K�<��C�o�F*���1
6��#�@.�{-��*�c�$=ފ%��6Fäl���p����w���}���s�^��� �Q�ޗ��xU�=X{5G��q�&^!-�5���!MH����!���:)��=���k��������P������P,
i!����d��~�����]�Z��'��N�be��1u.+پ��G�A!d��KP5tu�'��N���������5҈h��Hg�u�AԈ��"�S56Z��n����a+r��>�o�������8r��*VN{������Ɗħ
��*������- �T�bX��2V	$h��bI��N18�n�	�Ka����q�,^;v������_n�LQ���g�0K�ٛ���"�3o5ݕN�\��l�/���?.�hE�dX;fv�l,�Ґ7��G;�nl�sЋj6�Ñ
�Kh�����BQB�}w�Co���L�i�
��S��C�3��ހ�&q�G�;�K��JQ"�4\�W	� &���wp���bzB8c�9���dz���@��Q:��,M���g~.�����&qc��H��u!i��B�uD���=�#��[���T��ɹ�)N�ۖ34d��O�^��ZY���wd��_�5�|/�� ]V�ZZ�P�;�E��ZD�'?�餫&|����7�}���x�ܖz���KJ-ҊA׳���ʋc���o���V�N@
�ݝ�ׇ��<��W�x,��gz6���	0rP|��=�R�)���<������Ɉp���D�|�V�)�Q��u�\0{���^��=��ר���7ݷ�6�\;I/�I�g/�!w�󏨭�~����!؊S�L�t���P�������Y�y3�p.�z�o��i��sQ�m�іf�B�7s�A�z%�Y �mrީ��P�q�Tj��+�[y���|��=���pu�iFR�h�����	g]�La��y��5!zK(*�əl��*>�%|h�y4�p,�F�ʊ�#^Bݶ 
�Up2bF�'�u/�ɑ��v-p��H�:��/],�ȇ���B�P���x��+n�V�݀Yzv��n�� �Q�V:�ď��\��MV}$��J/��e�IM��0�H�j��_��b���H��Lk�ƘBDPύG�L5Ve�:�'1�-$��
zw����i@�Ǟ�N6ML�T��i`����Ɍ����z,��4��wf�����F����F!����cz��u#�F�qJ�a�����/o�����֤(�|�"ʗ�+��<��W�c�+�Z��!�l��%��u�2S~M���d
����lPW�Ma�lK���қ��:�LS-���_&�w�2(1�?�kX&3�^��ʦB{�t�&f��M辭V��F+��H�J�.[���o��n��	׮��C���gp]_,���"��6^)0���8.|�'��˭4�O��g�X���2?�՚�[˽@CW�lxe���5|܀��Y��Bc��/���&����b��,=����Y���ˍ�憉��ėMr6�\��X-f�6Ux��Cr�C\n�țY���Od��Ƌ�pZ�U|�r<~CQZhz���m��Zma:�E�*E�K�S*4���$\���g(�}h[��y<t��T��T�Z�1\�_8��_���.�A @E� u�}�A�%*n��k��d0�3�N�M��)(�*ݿJ�����`]�h-#2S*��p�i�Z��mT�� �5�ܸ��2��X\f�ҍ��B2�R*}�P9hb#w/s��3;�yh[�d=��?�����T�-h�,(�%5���Z{�mΏ��ms)�@�]�	�D��i ��Nz!�Z=��g4;>�r0F���<F�-Bfs�W�Fݦ̪
�ܛ��g��Cz ���Z�uP�= �J/Zx&]���K���.�����c	x{�i��	e�!:��"���~�Zb����-6�B�}�Ir���vт7���РHw�W��aX��V{���k/;_l�N��ve0^!�*�㢖Ι�hn���.s�M��y���� l��|��7�PR�/e�8(%�mE�v�;�?����s��yƒ��}�-�v�����l/������>��{��S��/#�-y����l�%�$��MFFk#`�d���x�L*uyc��@���� � �z��5�#[6رCσ%3�+3�?7Ua��3o+�ޥE�P'g�_�a�&<�ϚuSI�Ba/fc��i�&�\�@/u��餦���	k�҅A�����<�s,��q��"�A�6�4�|RW?�}�qۆ1�E/�@#c���_�V/�qBN��]"��3z�������|Hݎ~6��< tK��@3{�5��鵠�k�ʠ���`+l�����n"
5�`���5��Y��I�gz�T䀃��'
�R%�R�U��8����@�͠R�D�����5���.�=&x��E��ْ���>����R��Kء>"�c���@�OU]�g z��"���bX"�ޠ�����l���܉�1-q�?�I�b�Z�e�5���E���i�����iQ��Us�)]����x�}kU�$��A�i/��@��?dD�Z���U��OE���;`�~���r^�i@;N����|���OS:*�S���5{�+��U�7�ҳ��^qcQ�S�e��Z����"5��>'��D��!x�+����M;V~k���wR��b8��¬*ީ�I���)�-�)Ҍ�8W����P�vk"8G&S�!&�)v��*��k}a~�	�m�c=��P<�iƍ�����[/熯M�e�/����������
aE[��U�oݰ݈\o��O���jRi����1�?��҇�C�<#��N�L���Q-�ȭ}M߈«F�$�,��}W�"���xn�"�r�ZE�j�K*�o�8�!G͠KB֦��ډ06Jk�g�,}	)p�� ��a�xb?��[��7�u>�i����9���29��ɤ-gF������a�g~��D4ax]8;s�C�95�@:�
��@�[ѯ�A@4H�PC��r3g+�)�@��:��� \b�1x �
��[�@c��|��i@�6&��Ut� kl��P��)�HM���{b�f�(�`
�dQ�79d���	�<\����i@�"��r�Ҁ(��<���P����&�!W)=�~������M�p���oԚ��j�=�0B�w��;���H��?Ql_'�I>هVQ�hȵ	^�N(�Z���Nt}MprO\�}wR�#[9S:9�8 fЄ�8���B���h�y�j�O�	�C	�֊Z p��V��@n&�M���\�Fv�(1g��l��e1� =B!xV��	>��CPlU� ]�?����>x�����Y������:`��B�%��{�x��}k�"$�<��ZZ�ñ�.��ߡ��
.�U�q��
��^�����Z��P	9��~�-��5~J �/���U�}#$��1h��
�^�5`��&���{���I�׬�s��Y"���/�t}����n�!C�?����!��s����Ks,�mVhW#�4�7�ZЭH�R��5�:�υ�E�_<1������S�LP�8��-�4��x���|����nO#e�LEگǘ�
o!��8�<,��D
}�3����%� d3@�K����ٵ�'����:
Pg�`�:ݔK���3�$��F��Pu��?�}PH��TB���CG��o-���xHu
�Q)�1�c2�՞��dg=ߏ��|:��\[D>q��s�MP��vF���I��b�S�d/���qu��M��K��-��P��B	�D�=�M;W���.s^
��nV�R�\F<=n�i��&o�A�s)�7	�<�@������Dk7��&�vپ84o&����QB�e����}t�"&�ȯ���
�h�\mW4)���Y#�i��z=��4�]VR��0O^W��}I�i]� �:���5o6���p�����d���	X�PfW6Df�c̒8  e���Z��J��|fS���s:�4&��uAE�ń_o���qy_��"�d��񟋝�6�G�8VpJ\'���a�g6�:��Ӈ����G�R�=>����y��ӎ���M�룿�i�ޮ��l��ݨ�P�Ybk|%��G�2�J��ݽ�1��L������^\�N�y����)��@���N0V������#1�q�����1����!u���c�A�����T1C1qq�MCo�*��*��S}��w����1�@y�Ki�Lz���E9 ʷG&ϫ�<��J����&")MI<�6��-C�j b^���Y.����&h��Z_���40U�ⲏ�.�L���â/k������Ed�/{K= ܘ8�c��έ�g*D䌏��w�t�xXA�W�0����$���zG��c�^M=_��?䑇�Y] ���+&{^�J~��U����X�6}B�:8�Ϗ���ǿ%m�TqWr'� ��Sj�,�k���H�|�mP����i���u���;8>++���[Zg�KXG��<�c�A��i��P�Zi��1��@�v8�������<{��!��F9-��H��ǔ��\4�k��W�(fh��0z�q�<M�uV��8Ha�::�&)1��ܯkn���K��y�0���*Eh��a��7�cX_~����z��L�����3�<��~�.f�����罠��2�~ b�	��YQ���I2��K�J���`x"}�~@���43W �����{�"G�*v!�\+�)�K�d5�6�z���	��@E*G�a��*v���1��ýT^���L)�TU��8> ��Ut�F��]��\����#�e��Z�q>t�FE��_���1f�2),�����Y�Z�c����+tE!P�r�~l��Y3t�+�9��4+r����HV�#���L�������$`�V;;7�sS�n��y���L�>�̲�Gf%���(�E%fv ir>b��gO78�V5�auD�޳���%O��<:e���8��H��>DN�ǂ���0����ϫ�0h�o*�a�I�U��������և��Fv�a�Fy�G�g���	�$o�SQ�c6���Cڋ�ش���� ��1x��<�ԩ���y�2l���w\�dTgB`� ����{�E�UԳ��Y#��F�cL�l����miV�����B���./�K,�i�ٻ���='���MQ�d���mP��������g)��=}(qg*4�>�p�B)�@oѓ)^�ko@�/ ��_�b\ ���k�A�=��!�g�]�s_[?�
�6v�LB�jvr�Z�%�j�Z:$�t^�Fu��-�5�/Ԥ�+4!wr' �KPOX�|;����Q4r�Ty�ɑ��O'�W��Y�7�$���I�f�=��9�~�"��(H̽,��_���#�?X;w܀1S�kP���!��&�'��"��7R�������+2t����܎�L�8py�<��W"����HYe�J9��_�$8h�[���W��o���$�]���q�]����jf ��P,b0���d�!`޺a��\���V��c=Ȱ��]�y��,O��b���C�P�{��+UO�\�����/p(�����g�F��gf�n�m�8JZ�+(�rq����d�Y%�89��PO	p��݌���@�8�KӐA�IAϘy%��F�}|[a������'��:�(~$�㞷��A[��f:��<K��s�盶�4ʓvA�.D���z�/)���\�٧/�k~��l�/6(�I3H���B*\܊�g܏S�ѭ��9�)Ë0����^](�*�̛�$/��6s0r���ڨÈ�)#,�u2g�ʫ�c�O�ȕ_�H'AI�jY���/�����ʢ�h%���O�,��]P�U��؅��Z@�w)���F?�h+����C-����d�LҌt\Ų ��6���H�ʸ�����3����Q}�P��k�vB�������X�85��-��|<�A� �U+ ���$(��xC�
9�	�Y��<q(��w����%�̤uf�M��i�o��Q�=� �G����f��f��0ΒX�.n^�}�κ��
���C� ��ٮ`��ۂ��Zպ�m�qt红�j9"�'ܷ�U�E��D����=S,]t[�����n�;�T,;{vynE��s�.��CU7�M6���� k�b��~_�L�Z��75X~�=q~���2Mv"�9�gcu��5EID��2�6'�Y�~d���#D���6'o���n��^�+i�y�H9iUw"0�]�3�"�5�C�+!�Jz�7�f�U��>�3-�lxC���JdU�fO�w �2�����]V��8���pҩ���}��Bi%����>� R1� W{�x�-e�#�)Kʦ�G�÷�aR	pp�!N��F�e�}�MX"��X��=D�b�(��l�i�@��|:L�c�c�(v�~�Y �z��S�#w��؟y_h��ص�]rgI�uHT��;bP��$�P3���p�?��ȵ+S<��fR۲����!S�^s�;�-f޾(Q�M�*E���^d��	�xe��z�`��U��y��77C���d�F�#�̬�S��뢗[�n�(�Z38�q�M�`���-��k_Ċ&XChaM
�J���Η`�gVC9@�}y�s�{Eg!�Plq�#�;_c�+�?Z��/��]E��J%A0�~��P�q��Y!fQ��� ��kȹL�'�K5�up���0b�U�|�8u��5�2�z?��¿�`�m����v��d�|V��-�j��;�~V#��=zG�Y�.�F�d��y�/S��%Exb���NN��/C�&�|@��t���e>����shr�V��=��g�>��VT�)i����z�2\YW�e���;Rr*��WeA�Q�p٭�A�^�S������瞭���7i|����Bn+��{���(?��/�OZ1���c��i~���eo��A��wY-��#h-���t�ڋ�ɟ��ah��οR�p��T&$�b�S��ZA]c��TS�H��Xj���ϒ���F^������[LF���<�V?t,��f�*?zKO��\���(	��)�	��\�y�3H�~ьK���'��ҁ3�-i��c��OB9Ԑ#3������JV/gD�g�����&K��S	�������j�6o�ng���q4�|�� ����0�WXx���x+���-�E�=��ԗWτo�a�:�G2O����Z#�ť^�z6��I�yG�}?I�l���)%K-��C��8q�ĠX:�L:k��Y�X��v�z�2V�u�q�Θ� ��N�dOk��6:�x6�#J��blb��hl�� �u��b����䚛��(�+�7ßSo����<�W�
�����g�N�j��� �����`�J[^�]��yh�����Bo�
�������#SWJ�"5Yq�WC�f@�k� �n3�W�y��l;�N�Ev��|s=y��W�%�%����~[��@���gx�ph�ݓ �%������uW�#'�҈���H���Rt��S}�W�L���ny4�Q�� *+H�1�7}���&M�gّ\Pa�u\=��d�`�@&Ah����i��@�p`CXP]gφ�顊�[Z��&KӳC��}F�=����"	���M�pE�j*�]��Ӽ8�C���U�CW�ZJ;¤�~�]G�-[�6r�ؒ����--���bj�&�:� {1����*�o�&н���֕��)H��V���*�����㌕%�؜�(K�-ۀm��-�I��mPF'�����+�Y�R��{����ߛ,�fN�HF���/�K�0���s���AtK��h��A�:w�c�R�`�?�6ly'��H_�v"����OƩ��EBF��&.���p���.��@j�y��F�>@�룩N#ܢǔ��>�%���2�}��u��j����#�����~;��?n����Ԏ�R���5Ny�3�NM���U��jI�h��c�����V&����ӏe���� �nH�\Nיܶ[���pi% �Eh�f�F�0X�2̱�˝K�0CKee�>Q��цnmЎ|K!'�{�E!Dt���r�2���18I� �'�ޫ�'��1�58�&�C-O�s%�'W�EmC_/"~��T":����XN�Ͱd�:����y��I��`��D���`�����i;`ÿ��7ן�l�5Y5���o��kmH��7ܻ��g�+���+��d���X�!�?�SR���bO
5�Y3a��#bdo�_Tx�GV�5o��tv����`3�� 5��!Ɗ\u���/ܣ�s��"����n}u���J*�v�wiwvo䠮����:�U����\����e��J���O���u���V���St�dR^1����z�r��%�g��G�0!:c�'��?i2YxX@��_B�Cal5�a��p�S�'N��&�t�歬��O�8�����Q�t�5�6n?8l!�"b.��+e�H�WL���c������=�)T�y'ɢ!1@h�6�62Jǉ���q	j�r}�� ���Q��?������$#<�jD�^���r�YF�*J�$	�;=�m�v����ׂȈ�S���憼���F��隌�Vy���-U��(�ao$��ߓH��dԩ)H0ۭV�ܸ"�"}FO�9U�B����3���7RȢ̵�N��M'��Z7��<��s�����.�4�y}���&(��崸�J�G��/