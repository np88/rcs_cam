XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��@�����I�F]:�~��ϵ��H���5��$�[��u�lm^g�s� ����~[X�r�Np��������Y����)���k=��A��:̐n@*�']5U�i�d"*ѐlK�*�{���V$�j.����$q²�CPd$*������!S��k��Z�� ��8(X�O�+�
��im��G9K����Hb�y��կ�y�F k���V���}5'��1�xJ�	0��_=}�TהY�&]��� 9�9۪����ڷl�Zq���p]��Ot�hyF�衛D&�!��)�|���Oũ��^�,��/CҐZZA�h��Gz�?�|U�~��UW}�o.T-�"�C}�����B!A1�ײ����'�`&��Y����P��n0_,�X1T^����ѕ�l�/Z���$�I���1�>�+N�>�<I<$��e���b.H��� U"�b��,���zO�gD�C���eY���[�����s���V��eܰ3򘑿(�8��t��1�m���l����n\�T 	è�������2m��J��H������ �B�Zy��n�]{�
��%wO����*&�z�w�ܙ��@r����1��ׯkCB-�3�N�iZ�*sv��_��yQ�/5(/�5u��N$�,0�� \ٽ:q������"2K�l��GA��vGV5��ݲ�4"�7 ����ӳ��h�*�o��@:g;( {m��5䒑��ߠ�mo�疋W*����or�*�Ȱq	g��� �g��bXlxVHYEB    117a     710�{|��,?}�:�Ecn�:/1�K�LF������:���el���u�2��)������p4I��ttD� 	5��@�@�OK�n5e(�����亀���Yk�3�[�q8д��w��
��X�At���i,4sW�p��gv'wD���|���[��m��^�]k��gH�����c(i��Sm	n�,�Ím�7�S8��T���|��'eR M&�63�}N�b�m�t� �����ǗcF��=�6~4��
ؽ��|�p{S{�RZ$9I�����Q��q�X�p���a>�\��ͫw\�����=p�j�7���o�񐛈����P ��9ky�����y| Mn#���tKN�&Gn����;�Z�e�/s2f D���p����M�a���. �ϓ1'T�BX]�a�Z
�0;������:�}>tc�~|�	�?,2��Y>�.t��s0B�'��dV���ȶ�K�����$)k��z���n���(�'�S�A�ťz�s��D�<��
����a|�~x�~�e!�>� "���{�h������V�^B�v�*�fܥ��ع��'��I�kX�g�bD�$�%L��f�����n����J���C`����K�T�����3U�<����NX��[Z����M�dֆ�%e��O׏Zm��Z4<�׼�2@��qBL����y�Ь���� U�t��V:3ʹT���}�����}W�Ra��l��
���J���(�BkD̰TN��mHq����ͥP�� xR��e�K�#��*�����
������hsN�g��H@s`�Lg�[�ݱ��˓���Ѕk!k��BǱ3����X��T��oW�IQ����ڞ$��6�kG�ư��8W��Y�����0��\����
u�*
�.���,*��lS;���|��sH)��
���[4-:h����?:��D����h�9��û��^5
Dl�\�#X��:�i�錇	E�9����9 ����y��t$�������%ɽ�.���8<���F1iL^f!��c�uN�qV�5u7���L�V�j��me|{u�>��C]��x�Hq��N����$��r��\���|Ҧ�z�~-�{��0ya��J#3���[�u�W1B�IUO忹��cje��J�iE�(e4[��?��������&-gI6o���4 OV�cW
�yFy�C�GX�_K�#zQ^
�jǐ����\Ø��׊�>�d� �>�~u���(�0?�8��x`X��'�I���^�~e����J�P����e�70�`��'��֐���-��!B�d�_�+��O᮴���ţ��}CK�Y���6$���p��S!�@��N�����PG����g�V1��QђЪ��IɁ +��L����0�4���n�3�"dɒO,�~~�|ǂ�C��I�p�mqw���v�bq���,��տ*��`-��e�\0��U�s��=f��^�xv�p�PMi�>�n�Ļ�y�>e�	�-�	��Ș܇#,�D�f�\�I[s�cMS���̎��9��.r�����~���\�l��2t(�W�d�z�����:g<�F� E�����D�t������,�3L���_z��b��� !�i�MF��Ę}w6�J�]��PϚr?�
��B�E�5��3�
�Yg�+�2��$�d`�=T,Ay�5w���u��V!���J�J�L�]��u6�g(��C�f�a��BM�т�*3D���}u��;�]���S��%������g��.�!�