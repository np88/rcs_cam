XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��o]	U�꓃N�}/�Lw�r�6c�g���Z��J {_�[ƽ}��.�AJ�28w�}\9���z'd���n$��b���I��9�E�A��a ��������Ɖ��`����EN��5��V0�h$�P�ͬ�C���6R�y\)U��?���@��ೇ�ܺ�����q+�/�ae&c�<3s�N�f#g���wr������y�d]հ��ո�o]�3*�󕟵������KRx�2�9`�hxw�d
�k�y���8�2�(���ugfT�CUP�s	���)V$��E*d��#g���Nx��K�S�,��ǻ�Q�����a
��ߥ*�V�(�S�/���x��-���2{2�Q�A�Z@�RM�Q$¾��º�)q���Xw���yp�Z��N����BE��e�5)yfq����v���Yy�q�&��z�F����#��H��l��jO=Wϐ��R~����TK��$�xϴ\�$���
kR3w���)�����J�J��=�B�Q�|<J�1&��wy�c�Z�TB��s'OHc`K9D���,�;�E��K��|'o�����/a��*��1ǫ8�C�0k�y���++�,E�	]Qi��'Qm�c��P�q�4q��ut"�"�ͣK�w��Z}�k�0 }��K�����ή	�e.���M��QlQ�t�
!?&Yr�N��)��6���P�p{*�e��!�SCHkR�'"1����.G4��U��G	5��~�5�����a�)Z�'ᘦ��)n�+�0�E�XlxVHYEB    fa00    28c0^m�[�AN�`W�=���pD�w�\,��ʘ�<nG] |��|'z���z�(yLcB��Ο��x4�?d���U�D@?ɟ9���_ʺ��藫��K����A�	Mm���m�ֵ@c"�WF�݋;T�:y��R.O��8c!	�+��z�z�(B�M���6�!+~��-���[u�k�(�d��!���$���>.�`v951}s��4 �jD˴3���2��g��̅.�Y-b/ڃ���qo�/pZ�d2E�F/"`i`=P�W kd��=
�Nȭ�k�d��F!8V�lM�<G��#�g��Ç�S�Tn�_�J��D_��`�Z�J(���ߋ �P������~�M4n$O���drQ�d�Gjx'Ma%�r�u������q�ؒp���]���+�8㭟(t;\����gM��.��c��N��n��΃<�] 5D2O�j�̈���0�\�h˥>ڭ[����:�U���c��H1^s�W�ׂU��.�/�il����6�j�"=D��_���vEF���}��_~��4�cy������ٚͱl�M�0���Aك��c&�!boB��Q����i|�Hbd�����o)F�U�JG���7���a,���S�X�A��g��./����К�6�Ʈ�����OJ�aw�J�z�R�Z�z�ˊC0*�t}�al�����]�9M�dp��P���M�tv�Db{nÓ4�� �I��.�����X��Fx�fX�	��ΡjF��=�;�(�ko�뤷l�v�ۀK��Pis�vTGL��E�<QVF��Ǚ�.�Fr��Wx��-���l����B�
�Ï���'ݵ@�����mTJ!�v�%��qBtL��G�~)s��n�	�v���Z8O��H����4�HsqR�Y�n��
�����'�8�Z_��AN�RÄ~ț��g�y�����������Cb-~��"�G�y[/'o"L�2�<D��|���S=8�z��f�{^�B� ^�s�2Ʌ��U�`r�\�F��Ԛ8'�:�����d92gJ}��8^}�������ba��W��-a�ZS�!�y�Z�)1������(^f	�ճ=��Ш�־��� �c|�i�GoV���BIV�WH%�����;Ы|_���M΋�[�][{ z��'k[C�F����
���	Ĕ�3d�j���}c	�f�RڑZ��ơ�(���Z/��u��B�e�7�����ॐ�h?.r��F���I�1���T�����y�^���u��<��Iu>��v��"�?2vw��ye�����K���+�x�¡}hs�@\�H�M@@g��U.����!�ꊇJ��>��w�*�Xq���>��f�/7�φ����@��q��u����Y��ųf~��2#k�'�t�Pr7��o�}��h�]�ܿ���q �Y��n�mV�'�M3�-_�����id��&>�H��pT��*iؔ�7��j��M|pD�^
�4'��8��o�8�\)�,(�f�=�.D��k�Yպߋ��g2�B���vֱ�3�6PX�H�B*Us*r�quF�h�>]��I*f��^�h��c��o�&B�R�t�F���YAj���@�]T̻y��!xm]��8ט<��k��ф�}�W��2�jN�=�Yƨ�U*�yv?�1-	-$q2fS":�f�qƕ&dL��ٶ�S�Q�u>ŭ������	5�=G|8�,�<��E:DN�������;Qdc �4�;��r\X��;O�Üݾ�O�ɟ%N7�0�t��  ��LJ�q�P��!V�
 _�X_NL��}'��>SM].=�V0;ɍ�?	[U�n"O����|f���$��>�g}�m�����`%�Դ�;I?@Q2�.�ks�{o*�&Kn� �-,�F�!kup��0D��\>�����& OIn� �����Ş�2����IW�n�81O:��|��@R�'dn�_�U�����eZ�-�l$��[�����JX�]�g��|F�b7��޴U�ՉA!��9����	fjE��k)X��ۦ�-�8��\���u�zf\�-��!1�M0[�Kcب��h��Ґ$�����2�<�%��zk�f��@y��Qۖ������u-~��,='o�3*���^8�/[�[���殈�D�����cj�+�����K��^/���u:�N^<}�_'
y��%��J��6��>efᲘ*�!hȾK�׀���w_���g�H���~D�oyJ�Y6ǡ�Hdadgs����d,P�@�����c65�\M�#?6�r
�>^����V�хKC �A���0�{WuYē����Ғ���x�)��m���CD�
���0���ٔe�w�&�A����Do3@;@~dͲ�����Da+��36"�Ҳ���%���!Ӣ�[Vd�>�?�t�v����2�U��>���I�O�У���؉Y�(-��� \6Ƭ����n��ͿX�}��t�N#_���*�Um�z��հ�'$aC��������e0/�x�
�&߳��Y��r�atk��m�p���Fe)2X�������4�?�	7�D!�G���_;Lc���X�6 9�b���W.@8��8b&::�ݥ�=��NK���a�FQ�h�.��`	!G? ����Q瓃�L�=��1$:��
��I�=����(�.ݮ������1���^�U�~�aWzd` ���?�$C�j��J-g/N���ޅ#H�v��bI����I �-U���
V��:�ӵ'�^��5�I)��&���bGl��e+6� z0��a��w�1�9?w���@��q��M"� *��p$zm�.������A�`KWu�o�Ӹ��Y��j��}���=e��r󽟟��������^�Bp9�'��l^�Q����шb1w3�2m_C��3�{3Q�J�\�q+������!z��Â|_��/!��}�c�Aշ�gw�Mҥq%=����b�ܙV`>�;�nv�Ʈ�:�v��2"e4�Y�XO������)%4���%z��ٺ���z����	4^&�2��RL�>�������]���Q�N�߆���Sh�3�������}	:��HtA����AHԌ������6��!�R�Z�A�=��n��Z� ċ{��?�x��R�頻�%�3x��	`������ɏ�ccC��v�^�M?��`��x��g~e,�-?)��'��Y��}���w���ɑ0��r��1��:�%A��s�(Oh��ML�$�ה���LO�h䩈�ߒo�����i�/���Ә�\�	�ev�?�/���<�nP�������=�ǒ��T�	3�id�����X2�!��9����3�Й*�>#�5�@��-��kIC��Wf �M�CRŚ]�wJ����$��ܠ.���eZBƖAd;ǁ#OH}�x#�V����V��k �9�K��@\3�Lʧ��"��{�����
����\�߻�����Q��I��T�Ya�w��4��O>Zd��s��5U�,m��#��츿�Q�4����9�prl�|(-b�AY��3���U�@�[t��|~r<��o��S�8 ]�1�&����܆�s����������ç��a��1���:�:�˼;�o`���*9T:����+��TղA�m���m���BM�	M�o�IG���'�N�G8��BXX%�|oc>\۪�L��|3�[��+[���+���wOa|0s���A~�Hj+M�\n��V@1M1�99��<��|��
��8�5�-�Xk�E��y|C�H/-��A�<8h>~A��T���Z��D�c�Wmڛ6�������\�w �� �|��;(l���Y1ڟ�wI�
�i�e�|{�wS���c�:Y��O�Z� ��o�|#�s�Pւ
%�5=D����(�3�os�l�J	�Y�R��� o�4^#9́d�%�/�V8ꩌ�)�'��$���I� p���9�O�a���I�Wce�B~ېB��]���=�W%2�k�2��f)��st�!� 1@�*�\��u\w)���'�i��w�O�mB�7A�@������NX��Վ��t�'I$y�N��/�ǡ�Q���QhH�Z�_+� �Hj�Ke:����F`���NI��N�f���	�~�`a� �(�9�a�,���H��\5 f�� ����T#�fU)���l}��_b@hU�q��'ϙ�q��Q�;&Չu��Ř����k Z[aa0[�� ���Ω���R��`�~%kt�0�[�U�ys��ysVB�c��L�{_�z}�$>d�|���������j���f���e��O���(ң���r8�3��A�AY���t��o���T���d������o([3%��H���8�u����
W�x^����O�*jR>�X���E�4�0�>w�)M�f'Ԋ�(Uo�J'���8ץ,�&i��IEo�̼�A
��׳�/�9��8gdψ�o��_&b�Ou��G�jM
a����FySD�_���e<嗢�4m��ٸ"�����*�����U "���Ĭ/@KU�w׃d���/.�[.�G�?�>*Y������_�	�ݾ18N�fMIb�f:�$�H!�"z�73�wP˚������d�<�"�!p�LV0�F�G˛�؃����n���R��wDt�����r��sr��3K߱���.�ʿ��7�pK�U���@?��P�?5��F��S�+G����A3Z���{q\0C-�qx4�C�ݭ�o[��]� φ/�N�'�s�:�?���$'�ȱp�V�S�E(,�e�Ь[�����^s",3�������
�ɱ�t�}�e�F|�ͣN�\��MO̰��k�Гa�s�h3J�*����]$hj�&6�Qk�\��wб��i5��ŋ�n tMq�痁�z��r�B���]7 �����69�:p;��af���Z[�LiP�"԰j�DtE����o�bǢ�\҅0�,%��D��g ����
�7+��.��C~NGX9V�΂@��E)j/ұ�=B ���#ZV�D"�}�	V��9^�ۓ�9�\�R�~��9�(Y�F�5��O���N䰪d5h�N�[���
���������|�������
�l�7]�����п�~��+�y������:n������b���n��k"����d�X�Bu*n�8��f�s�ʷ��a&��.�O�G1vr�!j#$i�P�^#�$���;�l"�~��j���W)�HJ���#�+-��c��G�_��ծ�or�kNEQܤ����.c\]=���_���|ݰ����!�#�U0��y�|�c#�L�N�ac�(��@	(eDO@oq�U�!;upr��GNDjz��C�3[�F�\[�Qǁ	W�1yO�>�Y�g3�gZ���g2�c�d%�n��?b��Q�$�gy��Ĳ�ɵ4�T5��^`m�2��W��tJ��|ք~�&|��.���G���i��oTQQ��̙�y�&њ~�ڍ0�,Q�xI��??��o�}?�p̌�k�xG�lf�%E��& o������ Q��^u�	��uU�a���������K���1W��D���ٺ)������'�ɍ/�	�Ӿ��$� �p�F'wĚ~����� ���Y���B��B����x��O�۽E�U���>Y��@���:BisaA}}�[�l����c&&�&�@%��K�^���T�fhThB5�[֠��"�1�آ���]��vHb�2��k=��E��%��X�v�B9�$�`��;1�[�1mZ���""n˥��Q�'����ʹe"v�JN���T �K褜�5a"��V���ۡw�2�=���E����;{2��f	tYm�c��Q7e9�ap x�_ݚ� ��0��R0O����Ϙ���S.��_?v�C��"�Gǲ���C�،���E�3`^u0z�&��I4��8����2kL�+4f4�$�A_�7 B!0���4�P����v1L�5�&����Mu1���άFV����$.kg���!�P@L�B�c׈{�=%xZ�< �;Źh����hF�R9��L�k��k{�����n dGI���?��k7���<}Wx��K^X�݆���Y�-���^_C/+��K��l��A�y��5O�?,�3�p�%H<����������^Utꩡ�&V��g�w�m>�qu֒�0��.��Z�����W���0H���,��;?S�/��Ddx/P�irZ��u8�����,:��&�޾�Ak�t~��GsY�o2�i�*WʥgA��-�i��¼�P-�v��Kxs�~�%q	�8��4�s�8��!0�A�������ͤ�O2�ƹ���r�	�C.FL������a��\��7F����)��._E�j�"s��`/@�ڗj�w��>{�ձ��V>f9�Q��$!�n�0o�� �g^G��Z��Ui�� [�i_k<��)�T*w����6��Ň���kĳ/3���:����:0���C�\#+}j��ޕb��,�%�: �`��-J��m��*����\��d��a�M���I(����=w�c��B-c3GΝ��Њ�Q�[R�O�!%���������ˁ���)H�����^8Zq��!�NI�Z����=҉�F��_�z<J��-F�pfpK���
O�w��Z\90��^���f�!�n����%���{-SU�=��!���^,�z,�* W��IY:�TQ^8��,�V�)Q����|�n�ـ��Q[�ƉH^�K���)���L>��skn^��bΫ����?q�c�t��4�xi1k^�ﱪ�s.�i��g=�y���S�e��u�(�O9A$Dj�И'�í��Y���J:$!O�"�h��hB6�R=iq˾�J�H���N��j@pM|�"}�AG�I��oXToq�N�..m!�M���v|?4�x%�t{1��#E�f��"�-�L�0hW�0M7Җ�9a�.�[�>L5�C���B���s�g�
��Z���9o���p��j���O/M���1�l�[��k}&�DMN��ߨ������Q�?}Xu��L�;�3����9�7:f(�������
���gU�$˝�U8��<���;Ժ��D7���j��$�Q_���k��������d�Iv��(t���8Z��m\�"	hwp��G��Q����G7�J��x������`��}ghX�|��$��>�e�K���M��YXY�P�֝��@��.HjsU�7)t��_y���jt�q��k���� ��]��a���a��GyD�p@���� �݄ez����8��)�5J�@mU�Mg�=�Y�+|c��&Z�2ם[�`A�;��`c��*�f%�>�jV��W�cL�@}}���%T��{��9�ޫ������N^K�����^qލ@ր�lw����s�7����i�J�v��2{�h��Q^�i��"�sP]ޝyH�	����t�C�������E53l�=�(�zЛƚ;�:6�ж:���ۄ��Z]�H�*�}S�k�H=A���L�4E �2�E�Z�x+�K�������h!�k���C�|�%��������$q���D� J�=u�tF�Z?�q�O9K�3��$�k��q�f6�*M�S��h�m&���\��#����e��MPS���?��Q�;�����æ�)�8z�\	m	�0�Z5-�B�9^�B	p����87�u=�z�:�p6��t�e�v��R��|��ư�H�����PM����'|XSɊ��+����.��;�Y&6�貽���E�.���]���4��D$	u��ų�X?�홸Dd���)�����Qק��ۋOqh���}��1	��_��u�@�!�b ���=ɳ��� �ͰOri�{iH!���U�6�_<��9�2������>�%�%G�yte��ߞ:��Ո2�VW�J�Q5��oO9x��BpUA���z���-��U��-�'8�39;�Bq��%|��ٟ�#���!���mUԜ��l�K�qܮ��cgRZ��.�� @ )�$��iG8^<0ECn|�~��n����{�l
K	��8� (��9���q\>$t�A#�#����޺�p�;�Ҿ{dI(mŗ��^���] 
9<}^������?�x�g$�F3K�h�\�i�q�=�.������M�B���+B��>*9؈c'͊����b���C����a�cTu�T�������Ƿ�Hn\�A���IX��8�¶�
��u���1��T5��\�0�� ���ꤕ��Y1�AN�<H��|��ʹS�
�f\.<<����
f0��<��<�<FE�RL�[k��+h����{ᢏp	S%@��5������$;<
�
ckT
���ݝߟǬ�)x�4�o}��N��������Z��}l`�6��oC4'mƦ����٤U.����3&��y+X>�`�����6B�;_��A��f����8��؈��r� ��8p}	A��ͪ0�sm�B���S��u�!.�����n��Z�T�͍Akx��n������M�Z�滘��u��L��X�ϼw|�{w���]�=�f�Wzy3�q8ܕ�SLq�����ACd�,m��&���]v�� ����k����.ِ�%�o��"��
�V1��a##�/�x�5Y |b�x�/�HպC�E�"����:��?'?�(� I ��`Onw�Dͮ�i�A7m	l�El�Of܍�y챟�rG�P�c$�u������z���[�mx���,y�8ݎ|4�5
V\M=�&55ЦA�_�dg��v�ƒ���~J�?jWd��&�x����׮r����C�ԭ��c�M�t�v��|ȟ����K���j9��P[T����}8]��h��r߈��d�nF�q�n���k������+�z����q��.xx)�M;״�3@�PA]�'|�q1f"����id����N��?�5P/X�
uɫ�r&(1;;d]�Z���?V)��Jbnq����﬛�fj�z��"�Ėa��T1��s�k|1�sFa����|�l�dʗ�uz4���qVE����
9�V�Y����ŤX�ηПp�z�|rq~v��Y�����F�]�����#魪��0��\RZ*�ͬ����3`�����8��5���!����Ԭ�iy'��6r7�{�D~���;���#��u�1�\Q�6Ѭ�@-,#����^������oI�K��H_S���^t$�淃��13�y�������6�^J/C'+�W��Q�h=�QQ.�c+�($@�BF�`ö��F�1]���@��Nط�.��9-g.�&b���h�U�e/�x߾B�ըǏ�i��&ϓu\��GY�>���=0�aN���h����
u��DigSv᩼x��~�m�)v��̊g�J��B.�� z�T<Y��B��ᮭ7���pt��nx
6��<y����!��Ǉ�:�7h ��"��Y$`�������Lg�֩C�����^�i�o��~��u)P婘�����Q���L�X�qx��=�e���h��ey�[�oVs�W����n!�o��O#S7lP)��A�D
����30�:8����Qa\1=�V�&���O$>j/�u�VZ{�W<ڢ .~{����2=�[�uTl��ӆ�H��+US� �-c)!�h�Xp����xR�c_j蘧�;f����5��T*tKμr���=,��M��,�4�Lʪ�}�g��\��
E`�W����B���~0J��0���wLb�dwE8Ni���D�[.{�0@eZ�7P�X��	��L�1���g�E�����	ü�\D�[����V�,0��mdg+��t�+�zy��,�~���Gp���2���*����K��)?��Ld�wA�,#�B�r>���Kbǲ�׋S
�OWs�M��yF2ncxT5P&�^[�(>$�#!�v��Ӥ���Yn���K�JQ�e|�z��Nzl�x��K(�6��0C�����ߒ��\5L����[c4ER�Q��u�s�!-��˨cЏBฺtƟ�<����dUO�P4�GǑ�|~V������gf�}v�|�1��>����Z�2&�m�z+��{6�/�g�G�����]e�ٿ�^:94�8S�����1;]	 Eh����39Iɠ���?��z(u��,���8�I�P<�Dc�5�C�2��[n�������W����4��4��z�ϰ+}m	�&+nK/���o#����#26N�<-�D�9��=��~ި6�XlxVHYEB     896     280�ʭ����b���[�!�wy�Kn����Fz<W}��ET��� ����y��.r����Q��A�C���	�|��{!"e4�\�R����V���X�]��x7Օ+��H�9������iG�צ��K_��@�_\�/w�[���q��A�)��@�c�q�m>���
�%��
!UwzmϽQ��9�t�DI`V����zP�w�H��,\+�]�L�8A��š"c>��(�:V� �I6S6�i?�x�	qfO�+��B��ml��P�a���񤤟���
��^�7?N�fr��E��
�嵧|]��g�y2���.�#*�XQ�Gay,9X��˰F�ǀ���u�p��:dɉԩ�.�B��JQ�LbC��Wp'���R(��i���#�mU�,礸�rZ�X�A�U��=m��yH��A�����2`�˕��N�2������_-�[Z���8�k�m=!�{28�F��%&Y�O�
�:>$�� ��b=���{�����;��i���$��ۋ���^�3錬띕�|�Zo��R�mH��[�@�i�44�d��Q��HO`s@��̕�Au�f+R�w��1�]u�_�+���+�E�
���i����봑�HS�ol�+@�x���� ��*x����n��,�7