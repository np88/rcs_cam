XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��(a,���,,]���c��~��o6����O\}]�`Y@	s���W	�A+�˅���r�SmcᏇ��e"U�ejU��1��4���ғ�MI-}:u��T�ɾK2t��7��V=��[��&������lJ���;M:��kٚ�?'�����_X���_�����IҜsq7l�$��-�O�>���(W��m�8��I�
Y�B0����\���g�A �F#*�2�K����;r��	#XT��ft0a�E'z�b!3b�y_P�ɿ����փ�D�?j,*l�-��)�t#��9)�4����J�˯.������M�$�nm	�/[&Y�A�~⧮�����Ȃ�jHӝ�Wq޲�s_l�d]n�?�aZ�,
{y�M���a���ޭ�3��y��n�O��o#��7��&�����Ћ�|��-�={�/���p\3B�ƶ��a���h�Hlb�k���R�����Ê�v��S78E���N��/v31�U=�N����/=�K`�}�^Y�U�"���U?V��Qxĳ:��L:���O0*(9E��_�T�i�`�<��ax�#�;r��!���Xo��Z��R�W�U�נ���T��Tɽ�z�%��D-D ��t�����4�h����U)W,i� 2�f|M�sgq���{?�^��'J*JI_��H�*x��>��{��WG�$��c���@|J�D�`G���@�{�L�x��ۻ��S(���ޮ ɪ�'l��TU���i��y���'7oXlxVHYEB    33bb     c90
��p�(S4F7Z	Sm!h��v�����ݯ��˩��k�9U`' � 7�=3���1��B ���`��q�	�er�U��W'�Jk����⟃���;V���.V���8�A�D|-�������TO�ݑ�kp�~��9Hm��Z��rQ���R:h���cWDJ��g���v;l�#b�������_�ˌQ,��aN�6aY�P�l��,�������~��gK�D�*�el��Q{�DOJ�6m� �9Q%��А��ˤ=�T���dd�h�3�L��3z泬X�x6���邹�3ۘ��](r��v��L
XAC�F�]8غ����Ы>6��@f��pjT��&�O�m)ʭ�c,s�󵄐�sر���� +����1��}%]���+;���aj-ψ8� T���?���%�%䯗�HI^C�Z����y(IݿjV������-a��s_@ޅe���fx�Wv�D��:�fъ�l\�{}k����fF�n5Cjo�鵧���޾	�#�sH�Q�� ' ���5]�LWﶦ���o:��UZ���GnN;�������V:�M|ޝ0��98��a*`��`�tx]�I'��U����:��G�k���3�BX�>wS��7�5���֣z��j����^5�a����oy��T1ޚ+W�ߞ�6[\ϜQ����+]�If�e��D�K��hn�P� ����_��׈3��x���F�Μ�Z c.1f�m����>��X���@Y�q`�3�,�i�N��d,=%!:�w�����J��'�/Տ��U"���<���r:!`���T}j ��v �}��d!9[�5�ұ��-J8�����W���匲��?!�c���$��~M^���2\��Pq�B�aᰳ��>bP�ߤ�N��&���
C9���j\z@D\'�3`�p�~���f��K���@{���`��>Y'N�: 7���]� �.���\!r��:���4�)k��6�s�;�z��b�BX���]�YI���q��?J����*I�Ԓ@�(��M�_|wyw��f�}�J"�i! �4u��`<�!�w� ͬ�����{�ܫ校���/��/�u	H�Vg^�X�E _k-N%R���fQ/�}��z��%8_s��Ͷ`P.lJpH�}�6�Y�&Y�Xn�3�Jep6�OR3S��[hj+?��Nuove���#&���L��@�?��.�P��ͼ��J�V���'�~���@K����x�@}�/������Y2n��n	S�ȍ���}A����>[��uG��ns�H2e��˰�q*�������yؑW��p�����oFƕ~҇����
ʼyYV�H�}?U�u��Mn� }�ϝ�� E7��Zg.O��ҽ�Q �k~	��u�QiE��U�y��m�y��%π�����>�_f������M�oI\��4I�P3G�AV�Db���׭�+q�%Ǩ�=�I*t�:g\�R׵)N��W�]ڼ�������WWj-�N�o��pOfs�Ko�§����t�"w�JZ�B��1PCIt!�"�r�Ǽ^�M("�m�L��!�Qfb��_Kb�{�q�ퟤE���ʭ}�H���i��Q	!�͊�	�f�_ �;��)E�{����5G�cv�+��~:�K��@�'%�w���^"�y9�����|�ҧC���GT��P�ۮ�?j�4�Jvtn�3�Q�aʡ�M����t���"3s����� Z`3�n'�����A��2�kP,P�&@��{։��i �/����A�@����&���]�Ju�4��� P�m^��e����߹��-�;d��?��3��@�PjH'�tK�[j�>Tm��	f�"B'��$u�lW���H4��$D��fC�W�+�1rj�$�<m�qfy�n���#��ǅ|G�BY.�
Sd�ob��GM�A�ԧ~�S�`��d�J/P�	Rd�<MW a�d9�J
����Hyh&X l���+�J�DX���
�6�����4��Pogru�P<�L����`C��!8:T�jD��dA{��]9�*�T���kO\����^\����5A[�᮰��{�ݑ��	��7TDՏ�Y�k�B�
����Z������m���nҖ�^.Lf
��W�+c�Ѭ��x(��1��b���\��	0�@���|��M�d@�bOb��L��"��a�d��d;�{>�=j:�8u}�U$�v��S~�/�5*��&PAȑH���p��9��1Ɔ
]d�T��䠈�!AK��Z���m���&WMҠꄃb������#\�D�P��O�*�cd�7���D�����G�ȩ�����������k	)��|D8��r��{ݳ4d�1����3�˺H{�'�"k�g[0��9 OP�l������1ٖ�`��h1���\��
�v"�#<e����N�ѧ��Yy�sff�h}��s��������У��db`?ʠ@��J��0m�2{�W�[L5T���$Ϭ�̮mL���.0In���Y;	��8`���g�)g�"��*%��oɔ�FO]u>���g�`�orw_�o�h6�I�6�S��p�x6��<Cz� �c��{��8MH�F,�+aj
g��Tjd��ԥ�r�h_~��k&���I�֭���R�G�#�L��i�{���WG��{J��f�S-���̢hg��I�����
��.��q��N&���/8���bg4(��"�TX1�KO������.�*��m�M�B������W�`�ﻥ��%�d����m������*Y/��В9�75�aM6t���e�y)1Sڏ�:���Qj��s����]���-i��,F���w�t�	s�0F�Z�<6c*,���`�Z���sÑ/�W,��OݶF�Y��;�����R%
֌���-��Ad�U%�����\�ܞt���҃}1-1u�����[et�~��S��FZ�P�`��7-�S��z�� �=)�Q�6�6�==���)w��� ��{UH@I�޸jkfP7e��D���̬����ݿ�>
\	��dH�� x}�m	�i����S4gڢ�p$��b�;��P%��ʞ ��9E��`��4J�_P"�&���Z�Z�<�_ޡS�9�}X�u wN��6�g ar��y'��@����(f������P�#��	�0?r!�vNs4�� �E��V�ۈ9$�X�f�a�p8c