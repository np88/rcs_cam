XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����6�P���3� $p/w4G��u2�~�h����X)xf {䲴���4i��{o��+HP�Dv�$x���$�X��5�w>j�L��m�d����3��m�����M!�N�9�Id�s:ɕ�Xzd��,�[�t��oo�8���
�Ll��d��;��?��Ca* H侼�q�����s�>p��4�;�:XP��M��I{7�-����u>mA$B�U��-l���VOϺ��+9��Z�K��۩��C�h��:C�8cH!��l�T�F��M�O�A��O��]6oV)��qir4���B�?�@n\m�O�o���s�,\w%�
@�%���k��c����YwS�.j�uM�=k9��;]F-��A�@��t�MU}�6X�kyG����F
*t��?\�`-�_u�����>����<�N-����11�@�&|���xK턟����b��\��N!��I�
.�ߎX�z`TU^�)Hc���缚k���Z�zr|�J'ȭ�C{�t��"L�b�o4a�H`pyz(�����ħ_��̍5�gx�^�82A�@2��@��HP�r@$@��A���h*ϦZ�	zVEr�[˧�bsW�_��֣��W��:��S~�(}�a��59�;x���n}�{V~i3o�`_ur��R�Ї±2�<���r'����̾����aT��tʵ�%�+`���^�r��i|	���14}Z���+Ĩ���>���1X#�����bk0XlxVHYEB    4192     dd0�ٮ��WԪt����[w��qj��R�/���y�
Z[�:��)�b/�QM>�]k��?����}|`�r��C�q�]�#��=�S���0�&����πxV�z��Q7w�������� >^��}(e�bJJ4ӀB0��@xC#<�����_�������gàp},�E�خ\�2�:=� ���A5�t�M�ݠ
���-��0V0e�􈊪T�q"Z!CI��R[^w�u^��!ǪhI����:�3Z�[�w��J� �d�Y� 砍2�+Q�|�{�\i�g$<re�=�L.�m�5�y���M�2(���q�&�GD���7B���ǣ餦�@C�l,��hc�TD���#
!B����P�6)4�J������wTvg=S�cn|��
����\��{��EG�>�G�l�/f��o��H��r��
/�W���Ʉ|_���w�d�޷S��T;�	���\��v4�	�Z�0Þj��|��on�?���Y���oӳ������-T�X�3j�ퟔT"�������&ʗ�{ ���x�ғ���pK������aF��p(�3�P.��~�aI�.�YH�
��˻k���~��ٟzAk��z-V��7��3�Dך���k�d�e�������Eh#��@�t'%�A���>��N�,J-\�0�@�������{6R���V�q����g}�1?���*�m�NR�Y$���a�����s��L�;ݢ��� ����[�t��=}��+�����R�l] |-��0�%�^�G��A�T2�vj=�D�<	Rd3f�USȧ���`]���h�y�B�mp����/_���d�Y�#�>�reb�pB�P�^u�,�g�W~���a�&����B+^\X8�ݾ!t��U<���n��g�'�Y+y������W>�#A�J��5���=%�9�j�*��,�Z�W�?h�Ʀe��6iQ��~��p�����ڛ���=��mA�H:?f$©�{J��9��阯	���Ry�&�����&̪�����m��2F<���3O������#�# ו뛇�TN�����!f�����D�\,���2J6l��T_}�~�`���E4��uYՅe��Ԧ��Ŋ�2��hx3rx��3���f��H�z�J��L:7���OL�3��Mz�J�2A

����}��^�POC5	_���$D�5X�������Pm���5�غM�!u�T�����UN��E��1#��GT\����0� {]�0��'�'k��:�)s��e���͙?�,Qܺ�WT?3F��J�9c�]��<��x�Y>M���5�쾐g�lf��ܦ�mb
����CY���G���ɮ�y�M���1�W۝٫�ܗ:�g������yXF���7򋔯��P�Uy�9Z~^{��W5�S�2��m��[S�&��y��B���Lf�E�E\]Iҋ�Ӷ�О���B��+�s��g���GQ�M�q{���GO��t�M�b��	���&�N8���t�����b��%���N���:&��2S�����!�t���j����99Ж�g��lq���>!�"�3
�[Q�X�S��˳I�v`��E�&su@��uT	��c�/���Z��ON�2����Q%'�#���ygC�m	Ȉ�$�췃�߄Π�?��alB��_4΍�C����U#(�&���*�w;�(VyK��6���M�z��8TE���ް�=H�,`���⏝�� �G/�f��,�:k�lK�ܺ�X��.�F�q��hڜ�kD�/qp�(�P�iK8 wh��U�ޗqK��a�o~i�SPϏ�U�#?h�h��kj���(��m.��_TY["�_~7�W��[ZK����`��E�I>��gܵɈꡬ4�5�6N2��`
����,��3I�7��È+ʭ�P�9�~��̑�
��OM�5�b5J��m���T`�'#�����eb����Ӧ�]7e� _f� ����I_2��㖙��bk�%��h��4���擀�b�� )�9�� �����7��õ�ܚݚ�R�u�yo�x�Wz1�)aߏ�2BxKx��Ê��'��Z4�`<lB�]sF�qar�͢G��,9��q��n0��9O>]��[Q��"d��5����ܜƛ�y5�"��D��������l5�ީ ~%ow��G(}��S�7gT�V��m~&�[�X���Q�`�:b	��Y�ܾ6'»�b��k��<�5�����I�A>��&�-�F6�̑|�8��R.!?~�K���k�X����%�x�R3YK�J���X�Hkz�5'B��>K䎱��(Y&��YH���ɛ���4z��4Tk,�@@RZk���S�A�d��-�@aw��j���W�):K��Fl�u��j��o�PJ���q;li]�<�9$����[
%��'�t�wҞ��2�W�NOAx�m�t�g����̀������S:��m�U
UXh]�w�X[ �-]`�u��|<���2F=��ڊ'���� ��kBv�Fs�m|�TH��Y����s�~�a\%�Y��͠l^��y��EH��[M�g�Y��J{E�X��x��~�v@�U��4�`Ó7�?C;?�����f��oeH)Dc>ͪ�s�߭��4GCDc�_�ZNlJ4c�~C�j��;լOL�׮��� �����d�ڧC��<�Mq�O�""�v����- ��;�G�,L������
�g)1��Q��Y����:���$���]T�T�A�oI��dww��(��\t���'�<����7�M��SZ���Ma#a�q�lR�x�5�x���3��O�n}���2(4~��_#8e�G�B�|F����	����_e����lTR�d$WD�D�F^�UV��ve)���:��]B��^���}»��k^��Pv�y�f�}CNY��V���5�'�ԯ�ě����RI����{e�<���n�_B��C6�� �Z�}�����C��2G�L�(�Qv�|�}�\�\�X!� l.n��g�0�ȳ�t��{����0�q�H�K���Mꄣ����E�w�?�Ց�=1~�|���k��C��~��-�N���	�ۓ����k��f�p��LY�� >D%U�Gi��xq	T��:�b��bc���2�L���0.p[�ٸ��y�9��W���\9<���:�]�>1�O,�ׅ�ў�7�.�p}}�����2W�A��v������T��Ep"��jT�\�婴�q~�f<��#A�}nSg^q���W�S8��m����\��苒&�ͮ�\�u�Z����Ak�P߉�'���K�����[�!!_3�Y�y����b"]+yt�n`�q���F�j����Zm�8��J�}3��1fΞ@�qI�}T�ۏ���X\U����4 ���������5��Q~#l{���o��b.2sc����&�唔��X���	E��o����#�%yE%`9:�.e����c