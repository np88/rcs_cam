XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����@���{"x�,T1��y;!*�O�Uyi{�;�k�\]��g�S�tZR ��Oy_H�=�*u� �v����;��ZdFk6=��%�t��RgjE O����W_=�ySORH*��M�Ëz�ۀ~��4���cm�H��oĆ0x����ZjE� ��T�����@�����mX��, 7zW��L�;$����^���V� K:B6��?�Y����ǒN��KrC8f��ë�pU�j��v����?���ʷ�����>d���d��V��5"U{���q9�j����W�:YPZ�$�[4o�'�8�f����W-�L��'�+|5���~j$��{����v4%H���d���Wn���>�XR�O0$@�!�oݨ��SDH����eb1�������Eā8���ID4;�!O�����G"nc ��%���q�y��u���B?.�;����薣�1�2�?;�1ߋu�ׁ\*+��}�"I����$�bggO|%��H��`�i�^�5�m�,;��0����z�˓:�K��|4_/jw��v�S��c��Q�I4l����FD��m}���1p�e�_~�����jV1�ƈ糖K����΍.�Y��nNAvѻ"a���*`�Ӧ]��6�P���PƎ!�r��i�u! f��i�7~{Y����I��-�M}�Xe�PT�����mG�^���qg������8L?�.��<Ƶw6�dDHҟ ��x��؝b�����zs���2��rQh��#��%�b�	JcI��XlxVHYEB    130e     7a03D�>�������ãk�����I���;��"���LM�d�敌�A+����=��g�T���ݟը��S����훰^������=�X��1�J;�a��[^!cK�PWr͟���u@*����.������aU�6�o��m㈚Hu��(JTy�ᄝ�;�g0������u�b�A	���x��	��p�W �E�r�)��\�a���tZ��G��� }5�>�I�Z�;u�h?��A.ʇ���W�[@���<� ��`E]64�xc���U��o"�%` ����,��U;�W� �\���U���8ޖ��\n�W	��M�2V��I%��������&��h+
����gк^��M6�ip$(�yںh�J!�5\�sV/�1�$ڊ0=13 ��E�0��#����NӮ�ã�	ڈ���.e��+��^*E��T��|��#�Q��h�����
����l��:߭A� Aq`yl�RQ�A��lR]�9n�%��
uE�[߫}QJ���#A�%j>t�mt�a�gs�b�U!�I(?�a=�5l�Ud�A��8�0#���K�k����q���W�*������Xpj�:���ǻ##��Ѭ'�J,�EH1g��V�(>��S�2G���2hq������H�t���r�a/�yXH �e�`!���R��Q���,���:=e;Q�|��1 ��� .S���p7'xT�P�āa}���*�j�"Y�:Hc�����������J�=��`%倌��eHQ��W���y��Y[cz�ap���Y��i���c��\�t,��Y'���cCG-�Io��XT��$2�EK�b�=1T����N��!5����Q�*C�Q����R�v��	��>��L��ε\�a�����d�җJ�1m�a8��ϵ~��Hr,�xq�ꔢ�g`�ro���O7W�90(�\�aHŧ��ԁ�H�?wȠ������q+k���+	�h���\�!��r���Z���c=Tp|X��@:oh	ۼ!�L�\�0��tD���o�����H|*65��������\8�I��cWexh�eh�X�'y|�,�D�S�4�	�~&�H1���T�X���6����uVO<���/����6��]ǚe��,�{�O��Kep�Y5|�M'*����d�r�v�F\�Uhnf�ㅤxM�.��y!�e%t�ޅa��l�ΰ����tz��\CX��i����fiP�Ʀ��������-� �HG;�	3$r��h.-���_�C?��v��~����]�Cd��f�4�3S�Υͨd[�t�s"���R���3r���������3n2k�� �يP�&E��&�i���R��#�S���;pf�Q3����_z�����)Z-8�J�'`�Bքz]wF�A҆?��@��'�qd>����f�v�k$�c��\�Y%N�Et5"Y<f����.�2���'=(@�V��))e���w�̔S�m��s��
�Jf4��A�~�Ӓ=�S(�`9���W�zӾ�*�S40�}t#!m����� !u��/�)1;��R��n)�o��Y�MPie<9�n� ����l�������$������v3:�'�ٹ�`��~�� qw�a���#�����X7Î\�������y5�wK���)�Ͻr�~��6�w<Y�DMɼ	��.u�W�oPb�\���F���dCQ�zY[�$ޮQ@��o����G^v���Z����Gk��S9S� �����D�0���'"�ӂ�����A��K[wX}�ʿ��Jr�n��9Ո����J�[0X"�Ζ��p�Ծkw��Q�5)�UY�R���Wj1_��ڞ+�}�'O�*�A)5m��=�E$�n2�),)�0�Oڠ96����OZ�l
�Ҵ��G�B_`����WO}����)�J