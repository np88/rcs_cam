XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���v�}���X6-6�y�������ES=�%,�Gx�-;��" ����N��IĞ��~��;�F�qڨ�'�Rj�n����=���t�"������4XfW��@����EVg��L!�=)Q�hCQ(�����r�Q����+j����+�Ygp�	�|�,�q��l��h��F�ᇭX����)�-c�51�$T�P̐[m3����j��CK�ɽ�`3������1��� d��"�UjP&F~I+���l�����n)n/ z��Ll4R��$�Hք�P)\'�� Z;EQ��9?�z�Xq	��d	!�/��c�;:-����w ����uIA���DH�I[�O�����IِCaX�?ņ�K� �)�y��2��O�}婢�%�:��!)�u\lx��6fI�z�Us�ѷ����QvN�09>L�Я���cu/��܀�Y �l�#\����b_ �y4�F���sxJEf(�J��.���������}���)~T����?��8����ex{���)T� ��d�MQM�1ʜ���2+�^�m��k��c�����z�P]�+*�dLQ$DN�����o$H'�������4�ZK�f�F;��◅�;�A��*s�rf΂��O�Eg9����b_2L��Q7[�4�s|/@.�&]�l!���j;F#������JBƅnER����I�#��������m]rZ7Zz����̏BE���9���lp-�Q���*{jvc��P|���:fh�"XlxVHYEB    66ed    1670�J���{�����]�}|�%�2�D7M��E��Z>s��
�A�k�x}�뗽�Z(�(�p;`���p-�5��س��S����
lE�d��,�|8���b7F���ÿ��� Y�֜�N������y��_��8����\��!��0�H���w�_Ұ�x�2c�
0ؔ�O-���k��z2윖(�/�e�S���Z���LgK��1󚉼���W����rr0]��T��1O���O���l��>���kɤ��i������ �=�J���P��}�wX.���MN�X���5m��X�q�za-ę���I����Ux)rv��� 
6vP����y����.:[�8�
�G}�r��k���x�1D�
���Bc;(�r�(�!)Q�0cK}����F��>P�O��a�S!�ۅ
h��uh�OS\l;���%Ԑ[����T�Y��(
;���=y�H��@����F�p`f��5b��|B�C-䂹��d\u?�f�����J��ݕ��V��6�N^N@�Y��-�f<��j^:��\|nLS��} �$����FEG8�h�V"#�2x��,h�iqvs9��u�98�ך����K������I.�3E�y� ?��p�C}��u#'N�h�v��ūY�Y��W�L2�-fhB��Ԑ~�����D�R�����n�i���AN#�4�RP񤛰����Mw��ׅk���v� ̥���O��E,'�KK�p�?D��� �+J5ZA<�������|qm0��[各oe�|ړLb��}I��*Zη0FXF��\L�q���C�4@�'|��}u�v�,`vYZQU�Ic�w�"�\[�3�3�9q��o�G��:j��[�~2|@��o*�e�ar���6$�Uo�K�̮#ޘɘ��=ֆ��2���}�^	t��l�wS#2��.�����"UA6᜔�g�-��i᠖��^`G;B#\e�{g��C���w{ԉ��O�vV�H��x��_�Vp�_9w��͸�\}���6	�w��2�T=�
�e�	��w[dg�wmb���3r�*�SpNՖ`e>GXT�}���X!�)��C^R_k�U��g�WBZK�pCI�����:�#f��<Z��Ｙ�i�4�#���o�cz���'c�U~�2��e�>i�MSO��o�&�/D�t�qo���{i]7��S�]K�'h��U�p-������<ߊ*���ѱ6O5��7��+a'������*��|�� ,n������9����:��(Qs�F̐/+�&���[�7��h�
�z��NԄ��ND��o>��,�Gm�H���R>xx��Ssq3������6�.bp��,��фf�R�����f��H\HP�#�/0E���d��dy���=����j����7��`���zoE�R��*�9~깤>��z�D�-�?В����)�{8hػ\o[Em�+4�v�
�BfU�;z�\	K�<G����S]n�W�d6����Y�@଩�2��f�"Ą�v�rŵ�΄���sm>�Z���5�vͽ�G_4#��rš���f�p�����V�eG�;m��/����q|�gkf]�F�(�h���x���ǃ5Q�M��}@�0 OA� �U�r�O���XK.yO��!q@G��1܋��ԅB�I�A��8���������u8ɲ��ܚ"�4���C�`�����rtN �i������%2�iZ���=>(���p�)���&ȕ��C^ }�\k>C�V����hJ8Rq�f��dʃ���p�/x�nf��Ѳ~����߇Dh���#���"60ӣ7Y[�\�1���_��y`8$�ꖄ�=�6�e�E��Ӣ�Yeկ�XX�-D0yV�6���m�{���=q��RDc�&W���c��W6��ХO�uFN�e�'j\����4�*�O�,������^�:O[c��e��++��d-|�i~��bT�M(��JO��ץ��pvÍ$}�b<(���V1y�U3y��=)��ŔJm��JE���W��람g��Ol9^%h���Z"
�_���F�����9�������TEq�#I)U�l����:>G��ņ��؊^�6��%�"�]�?6��jԀ$�������Sc����IhQ%m:R��Cٴx����*Lê���g����d-�!;Ŗ����)�nB�Ð���y���w������q V����sjVG���� �
4�Σ<w�&a�]l�
�r��1�n��c2��:{�5�4�p �=h�ũ���-�9$W�����қ�TϽ����	� �ܧ�W�y�������]A
��t��Uz��"r"��5�g�?����p�0:\��.�5�$Ϻ�w 4�区cj1�����m�4u�p�N��pYT��&Ob�s>����iS��5�NX��l �|���W]>A\}X�ד��[[��k�%����Q�[��$��������V�-�t������9��A6^U�8�
���>gUu����$�gP�J;�}�
�ZkE`�:����1���LǮ���Es�"���K��:�s��E�!��J2�4�ge��?�h�k���O�`�7��T�ui�I��`�Ljg*�"nј�S9v����)Y��1OwC�oUal�D�^a�O�k���u�g�6&�����Ҧ�v&ұk��XW���W$|��� �A�����I#+� ��=]N:�iA��p[����\X�rAp����k�pg�m�H�������x-y�}�-����5n� 
{��B�{�G���Ĕ�o�'Է�L?=cs&����"�]A�e�X��wg�u�&�9��S����0{,���� ��/�=���A϶�3�H�q=���w0c+�����Lj�1Z�fe�/�u-�.�5O�����&/˅C�Ӕ9Ŝʘ��Z��f�Eݽ-P�E���EP��}���������&25�,��l�������ۀzElK�ʕ����.O�B_��No�%��3.*��iW�3"���b&KK�z����t�:W2�D��u?!"���j�k����筲=�1||�I�ז�
	ưՖ&o�:�T��W�|��^>��ȼQ_	��������_P7!`�ְ���x*��<c~Ԍ�K��ob�����7vB3��'�����Z��cm�����@v��0���p����ቇwf,P�]zL �M�:�rԞg�܀Q|L{���s�\���/��(�n)>Q~g8t\�9�9���
l��	r0b�N��	���R�O`�-!�pҗ��#泙}�e��*���Z���RXP-�����&��!�\cf�2iQj����~��_�Sf��6��^ݏ��E��=�X��7w��2	�����&.;���K֥�uNk��_�;����#_e<�(�&��2�G��ؓr�G��Ǳ�*CDR��á���!w}����rt�{��MLL-uܨ�k�I �$�T����l��н|��6�>��%*"I3����D�K?P�[��ys��}�Q���-)d`�ub��*����/�.�#ky���Z��QqWmcRD8���ւ���Z���_qYxq�$GMK=��.�'$	\�_���"��*Z-�nͩd�By���]ڵ��r��9�1��o�o��E
T1w�8�P�rP�|��.��-�3@"�Xe�P+P �������sR*�jY��(�G�'����)��\yz�ݍ�͑�^q2A�/C��@]�gM�{����KiY��Y��̠!��O�{������u�C�Q ԗ��RCP'���&m	l@�q�����8f��!�J�`#.S���ȶ+��X%����6��#��¸���1F���Õ�8��%:�� ��m�i��〹���N�1����N9nӧOs6<��FI�ִo��U���rފ����$�Y�#M0"k[������j�3������|E��I�m櫪�H���B!��h
&�t�:#�O1ܪ��P.0��M�S��"���h�J'S`�o<�?�/?����u������� w�S��%Ɣ�w\/��(���Ѱ��&O�k���n�6�k�P:E�ˑ&�-/l!^XԻ���H�g�i<Y�'\8�g+��dp�{ǉ�2�֛�U��;�w�4��ln=�֦�/=�A%I~��ؕ��*��e�O���+��u�P]ۋ�4��T3T�k�=U�X
EoI(�+�p������$���J�9�枊�K1���[E��]3����)ݱ+͉��	��E�+�>�p:th�X$ώ�>��O�"�n����iUH��%b���0��{�۷E(�AZl�az�C��I�l'�艋�=.a���b�����}�C��9Q,���-�P󗴦f�=�N�D;l��Yb��-"q#�k<&�W�nL��|&V
�D��������~5�)�@�],����w��Io��v�ڏ��~umi���g(�ѮmI�S���i�16��PƉ�ϋn^��C�'?j��ws�5U7��j��YB�F�ߺ-�h�\YZl����&�*ә��k<Q�~�~����f��h����ɘ�(���\V�d7{B�*�x�Ȫ5��4��(Ъ�H�x�|�J~�MV�Zѩ���0Yr�p�� Is��m��jрF���>
!!��~�A�j��nz�:H�߉�<���~�"~�C��<KV�����:�{BS;���E��A�tdͰ�T/��pN廬��v_����J������?���$Br��ŕ= ��$�Rp\��
�(�QKG>A"s�4���z�G��JYj�4�ɟ�ذh۩�b��ſ��<{�4�w�5��@[br�`.R�����>Ր=�>�wo����CAߥ��	4WV)�[LQ�˪1xuz`������g��aR���X���4͝k輅f/�"tc��@]��EX����.u8"j.eu�Q�k��R.��e�������l�	����Ǚ����S��+U~����@��{�}��9[�>�&�f�>u*�d|�W�D��D�e�Ɗ�T�(�ێ*�uV䈒��3a�uO�2�5�5ُ�LN��rn����N�^B3�D��L�ŝz~����QÚ�T�6�:�����M���(�+�p���$�k�}c�9���	��.��m�x��k�P�$���u���S�:�Ƒ��_]/�0����C>��'[����ė�/�tX]�N�3��0/�MA�ɕ���w�����y K�o�7g���9�0�%����S�	�t�J��Y���q�����ow�6�9�7B��o?�9�a��i_X��T1$X0-� ���0�Bh=^#�m�th�6A�ګj�V�����'���b�K~#��7
����b�z���!�'�I����}���r�qŅē{7 G8����XG��� 6��Z��e�7���%�Q,v�"�������=��5ĻU$i��qcCL�!6sO�E�ĵ���F� �u7�����:���[�0�W�A{SX�58`%W4j�lX�s�v �:�����Ue�p�jU�����\�>%��GHu���%���ѬFEZڞh����w�q�m�-n��9n1M�����;6��Zh�"cS�nH��B��