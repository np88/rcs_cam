XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��z�Fi�,"x��y��r�������^uء$ı�{��J��.	)�K��\X-'~2ڝ�2���τZ:���)�6 &t�<�Ym�����g�	�B��VU=���>� ��;b���{'",s�%��4T��/L�X�8���'�x����U��-!Ar�v�$�ѳ���=i���x6)�2�+�"Ve���Y�w��Y�E/�4j�_�����-��6�2���l�p��`�0i�X��J"=�,<6�z �s�	u���Ѵm ��^��]������̓�xH�c�zFFY�F#�Ly֢�Uo�w[��z���Nr��9��'��*�R�f��E������Ioo;��w�8�����ˈ[��g�����}�&�P��>9rz
�������'� ���V0Z�c����%���\�>ULZH��h(7�։p�mᴬ�Y+��S�٥��W��r��4���%h�E��t'�L���l�=Z�a�=W�댊��ث���#s�P^���!!|%DE<��j��lK�p��{�|O�����l�E3�E3g�z@N���r�A|uB�u����Hj�y! el�sљ���V�o	�)qk�Ȳ�c�=����(�a@�I���<=�/Y�%����`EH_��5�l�O�ܠ	Hru��9�+`���$ptB �1�2���L��t��>M �8TcSS$�N��qU��E�fĤ�T�|���,j����E<��"拪QǠN��w���l��LB�XlxVHYEB    2a4d     c10����fy7�Rـ�=3���V��O���V���$\"�D���~�1�U���D�Qjd���#ĊMƥ$�Y���Vg��b^�$���y�qF>9?7F�0��CiC�Ͼ�
\��n��+��F=<�I&�Hn�wM��5v�ѰK�a��q(<�m#V_��@S��6i��1hu���%�{�B֏O��L7Ah��Mn<r���$~�I<i���0�@K�a� Cy���05�/%����~x����2(,������S�ä�`�[�19e`�N;��8��	a�r�@+w�df��4��{��|H�	��T��7�X[�Q ���e�Vϧ����=�HO4�z0?4�rj�<��s��i*�=4E�6X vqU3��m�	������%���b�^�\���,8,rK.s��R��'�#:0_ȫ�����޿��׷H}��Y���ю�/�j!n&���C�X ��s؊�A��#qV��`Kw�TDNG�Z�q�F4v��d��>ԑ�4���ߊ�8h�;P�q����AE��yP/�7X�d<�v������@��!CG�e�H�1�nm�nMQV� \N��� W���� H���������rŮ,v�q?��T F1k����+�ɽ`&�2w\zoٕ;��~o9���BY +�5�O����4=����-�ȥ3��AR�1�ŕ�	Ǜt��LL�zY���l�}1{%գJS��@��lc)�L�| ���)N�X��6��_���i�/�S�j'P^N>�⏞�[�j �oc��m?�+��N�LU��G�nRn'����A�o�t�vO���1����p����u@9BeR2ƮV�m>��8��c7F���S�p{�E�1�4j�z�>ur�J�u��&OL�F�C�Vy�T�f&��"?. Wv�7�Wi5�bU���6��D�s��E�?�� :ڵ�����ݸ����c�ݯ�%{��U�T�rt�s5Y.7��w��v��[9P�G� �P=pp���:S��b���qǋg��P8�ˊ�ly�8ͫjOO�f�mL5)�����*m��� �Iq��#��d�8k�}�ݎY� ���ܤ�i{־I�S2�'��nv��mͽ_ ��w����n5�a5r����Z ��5^�U��K����ިB�:ج+;��c�aP�{�� ����g̶7]�G	�D�:Jy�9nV5��q$>�ɔ�Ts�9�^KS�o�����n��w�۝����Z�ݑh"ը�ߐlg:|����Ͼ�u?�Q�'�WaZ1F��Yē��i�[�o�r-�'[���x��P���h_��]�^񢉡k*֎���n{��*�˞�0��AK�[6��C2�� 1���ɊU$�ٖǈ�%ֿd�q�6L{��j����m?q�c+�R��N�y�=~�|����ce�T�jhV#�q�%�q�Қ&��� �e��=v>��r�N{J����h�J"�B����9�<����]a�.��gXMs*�B�����?T����v���#�)�7���{�����n5O��p7M�S'j�=N���b��k�ז��cP{��8~�
���*��[;�ki�O!�[��m��'�:(�-��j�����J��l�J燎0��^���3N��U���3s���:'}��X9�H� m,�=��>7�{�;	���u�0�̸�	�f��GN�լGp{������N�%��K�>o/ׅNO$�t�8�J��h�3������p��[�f�^� @��Q��זX=�eV����Q�e$瑆�H[�����A�i�m��rbV������ZP$�0��_��Sܮ�m� �^+|���;���؊��<�3����ңV��*��P�Οж��T�$t��G<�q�X ���$9d�Oc�Տ�3�J�I�C�y���������K_�m��<��XKcDf���=����fc=���\�ck�ֿ���.��v��W����e n�Ҷa�Z�^#�G� ����ě���͖�٪���ųH�ԁQ���;bUk�m�}D]ɐp�����2����]�"�i/�'�j��Wt�Z��hc�+WlLf���q����}N�[n�[��=0Gؾ`����
�Md;�m��H�>Gxq�h}�!�|�U�S>B��Y\�SN���|-�ְ$�O�҈R�!;	>]|�?�B�VBr�r��6�?#H4S�4�Y֐4��R��U:<�����������ϑM���*��**,�[�x��7}�ӭLa�P_���a�{��|w vNK�f�(}&���Q�r��e���S54ʒ�[[yM8u�¾E"x�$g�	wb[<Tǣ>m�D��JS7�T�d�I蜌��N�^� �c�u��]���bv�~-�
.>�˽���������%x.�_���ҝ�����pC���?�%߅}�3����s�-�$�l!G��*ؗއ)���/�����A�C�/�.���)�(��Xݾ��#���\Ba�_���/��}�X�w�C�|��H������!�'�!Ζ��&�ç�Qd�-Ԣ�V��[�g����n�+�<)P	��dD1�/�N]��eb��1��S
����с���AaJCH�P�6�
�n����x}r	���8�݊W��f��� P�f�v��$�s�9����\0sif�[��5�����Id̶�qQ\�hՏQ�lM%���*� '=I�d�����j	  K�e6��5�i63A��l�&�L,A6��-@�y�T;���[AS%X����$d���_�*,'��x�ϴ>vjM��160a�+�S�E�X�3�f(Ŵn��o���;M����ܨ�byvR��!�&" ��ZHI���������W���q��l@��F�8&c��L_����Q�lG�����L@]��e+7���BPc
���p=�[TB/K����K�h+[;�>0�d�r~���o�m�>��0�ʫ�^�q�y��Ӫ�#�����68)'�����6�$GÚ�n�B��0X�8���g'��U9��t���