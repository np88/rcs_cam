XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��i��B�mf���N@}�L�L�3d%���e ���ބ�ׅ�����h�
�o����.��)Pn��2���i�s��]ƂVy�-��-h���9�N�a�TZ^�a8���t�c] �~5U�=aB[�Q�k����"���=����M�F��%?䤠-+p~;�/�?j�E�~���]@��v����گv�x��i�=NOh�瑠N��d�͜|kvaG�F��
���n�߃��Ɏ�A؜��Ɩx���C�&�^y�eK�[���r^�����,<m��SF?K��5��`�#d4.|@ǹ�G�����B��Cіկa���@��y�
^/�OJB�5��¹d�������+ >[P��>�DI�]�1έT�hˋN� Y��ᶊ�����CBε�����Tv���t��3Ya���7^�Xc8�iA�UX=���a��G�_&�b�����d��R�e#�@b�[	�=N�y��h���Vo�%̕'W�ޕ�΋�~�*�!��{!��!cc8�w�;N���D��).�Ga���>���խ\K�_t��K�p-��o�����Ů��gFGFJ��L��Ҿ�o���LC�'|q��o�����#I<��`�w���9�ྲ�@rc04@��ڨ�@6��uP���A-P�l+�����r`�:~Y�du�%wI��l�U4�Kg���ˤ��{�d�;x�BC|�;��A��n\je�'� *�xtԩ"+���e(;�R��-D"uXlxVHYEB    6417    1280ۡp0E�v4���i�S�v󹞓C�dk03�W��Ut�^`Â[���eb��s�8Z�2ߦ�����hFץ�����IS�.xý��l�p�t�m(��;zR����x0���rcfu��'�V>�v��������Sͪo��`�1�6*�|�n���+p�EZO���r�O�ĊU��n#�7O�񷤗kM��[f�ط[�G�¢OmWe��E��;2��םJj�b�C��hV�����	!g�2�|q@���oF��¥�U���i��o��	C�B�
�h��׆�j��sbt���ޔ��
�.�h���$܇�+��l����wĞ��^�]$��ݨNl�5�x�ٗ�F�zb��2c|�PF}��~L�_�h���~���I$��,�����sh��K�'(�`�GgK��K�����J+-��brT!�^��=��z��&���y��H��������d���j8nH���P�� ���!�v5opҳb.h��Wf�|��B��,��Y�4y��h��"iڶ�qXe�!�ه��s���4��j3�<����akm_%o��<�q*|�w�I�p,���=���T\�H�(ՠ~��<0�WfY���n�k�̖�S^ϭ����E���z�#��ӽ�`���K�Y�)���k���&,�.kWɴu�4`ֺi��%,���q=��oU Z��ox8�-�a�?�LĔ3��l�;7�̃e!G"�Y��(
���v��������?�@w�8�������h�1��Ԥ�ԉe@|�h��I�a�����c�z���,'�kz����[@�����_`A�T���X����xz��V�aC:�z�)�L ;R<� �ؤ���-܊�.bB]ve����ggp�3�y�l�1k�]봵���d}
�;DP���|~"� hK4�I=�3ˆb��R�.P0C޿�W%�o(���o���2jj��4�'q:�x{�`G��?4���Q�A�A~�;&�K�h)y�
�}��RԎ��gI�%�:dx�"�#T�Ԡ��ApWH
>�K@S��}��$9ft�ysv�=��?ui�OhFۢ��۰�f�P[Z�z�"U6�=�#�u���(��</�c��#���!���iK�x��)�I��M�Y~��5�*�p"bi�j�A��{׆�@}?�C�Rf}R�K|�����f
�
�Ho>Xߧ����Yi�4#��$��&�!BA�aL���Ӷ̎j�"gJ�����$0���ˇ�s��pP�9*~�nU�����M��E�O�9�i��g�p�ꮐ��X�-_������ҭ�]��Z_ǭd`51Ŧ���H�\�T2���36�}_W8U�㉐K^.�I�ݰ/ذ7�=�r���{ˊW\:y�l�����ո����M�=N6�'�z13���wh�߈��N���T�I��-�+��!�Ӟ`@��j�T��fZ���~�"SE��f�r�ܟ�����kh
� �3�c�C��3a�%�~}�k�ڬ���x��,ܪ4J=��Šs/{߷};�
�����;�hK�D-_��z���w�O��N̬�_�u�ڱ��
�t���
�<���s�����G�5!7���MN�ᆶ��g��<e���DƴJ/1���7h������+dW�}�ߜO�;��/M��j�!�-���"�#�,arao�s��ݘ���4���Ru@T�F��)��N)=�kW�YD�ڛ;����j5P����K"�&tW�����+�0#^x�k�^�y��t[����k��������)UG����\��U����3�y�<�q7���*��(����tV���pg���a�veބ���ޫ����*t�XL���ÁG�ͧj�ڶ��`�G{�>��RZ����`�@Rͭ���>��Wx�lڃh�
��SL����G�Tʹ���U+mÀ�4L;���A'^�r���M!˝�ٷ6Xf�˫�c+���z��Bwm��b��*�=�:� �$��4���5[�����J?V��P1r9~��bxa?�*&l6��s���pR���x��W�|�-2g��g.۟l��TY�������j	Ļ*�9�#Yض7����]����A	?���.�Ѕl*��f2�k�:�` 7���)-f�,�Y��8j�'�#�}�l���u֮4(�L��Wr��*k8كS�^<���nwsZ�$�<��Tl"��bԍ���\��['�`�W�F�����6�s���1�I���XV�C��B��7#�G�R�m�PK�Ј��7W!6?Df���A��ًc�3rCSU|����'0J��-A���O�&��N�P�c��7�qL�F�,ԡ�d9Y����&��Z���Y���b!���A~,C�{'��׮�B�"��y 
�v���H�?#pc����r^A�{��urR�4n�H��v��.ٛ����53���b1��9/E�g�Z�Of/��*W0R -)��O:,�r͢�����Q�㰳+��G�����g�����q-il�Vh�h@��p8���'��}�A o���_Ǿ��]{����|�v!u�5+g�,2��@k{~�x�5������^Th|#�:��|�+����X7�ŗ���CULTb<��HȏM�8�3��LR�r�D�$���*���^H�t���=�s�$�3H���mܸ��sqw2��Q ���4�:ˉIE���D�7�Y�0�2���τI�Ak��x�E{g�d����uD,��Vo���2hL�U�YN7�c����V�"z2�h�C	GCN�s=E���6����^7l����<$l9Ӳ~���:�o�	<��Cb��$A�,O����aSA-�~��V[S�TZl�E�WE lXB%�7<���w_�Ȟe��M(���<�R�\"�]���	,�G)� z�a-���p�Ӭ컅cAr�yh�DVT
w3؊&١ץ���H|k�|���O�R�U�/�vi=^m*�3WH�w�ڟ9h�iH`��3D�oV �(o�'���m���	L���j �nhN��
caȃbI�u 7�tx��3�x9�}�z�����j�]n����layO<p�����t�p�"��Ր|�"��;}_m��=�Z�@w�_�|P ���c�6��,���͙��J�P�"C�0�wm'��,F��9}�,l��6 [������:�?��H�Y��v5|W�Y{o���������O1��J��h0�]!PL��*��6�t��
R�:�V��A0�f�<�v
��Ш$��/j����D_N�z�*��$�W�ƐKW<~�(whbi`P�~]��^/��Y`9��*rDx����B&x��Y�$�=�$o
�}z��1?�<�R��v��0'���ح�K�b�U66���p�\��9�1�zA�j�W%/S�� �u��f�(f,F>��Z�&Hd*a��:]N��p�?2�uVwD�a�[\T�T�7/�a/|0��%/��J1�����.�g۞X�/�B
~���hag�ķ���:�%-�J���h"�c��ޑ䐤���ٍ�x���l�/��J�b��SV2�`��2�F�p��oZ�cƘ:l[�|�v%�����Xx���-i�v�|Ѧ�cK�L~,.ʟ���ˆ��^Y�v����&���������%%�'�_n��`�y���l�9�~�L��� F%� �҈�雬>e���Q��R�uԇ[����2d������vc�=Þ��#������`�ķ
�3�dq2�S��	A�F^cyI�½
�<PA���hIξ�U� i�/���́������Cf㦼	��<���d��Ķ��������M�4,�4<=��s�j��ry�*��f����H
�q:�����9��Ÿ폰}k����:9�^ON�$�UB���&!_VVxD�H�/�v�Q5��q8�܈�AP�=���Oc�Qǡ��1���O<H}	�����睘h�nI`@ y��AH�$������~�n`�P͝BN�OF�l��*�(Ʌ�`���{�!����G&�����JL�����6(�	4�������qUϘF�i���]4lv]gF�e�閡����c_n�cTI�b$Q�S*�.� �6��Y�h a�c?7P�7?��(��`�%X�O�4$ކ�"��R�������[f�M^K"bz��&�l�0��4�|�)�I���,�x�\u�I�#m��vW�$C����EP�L0It�.R1�K�A�I�-�ڶw׭�� j0=���'u5��ڌ�]�{)?j/~ӕ�oK:���ٮ���+fU5m�,Co ~�*{�O�o��7�*&�H3��-�#IT�Z�}9�6�v}&�%Hq�^���Iv��y�
���W��]��>�;x0�V9?���`�<���8��(z�j��	X:�u�U�o �=B�&����WDɬ�oJ:����y���+��&֭�o���']�|u�خ�{8͹ܯ����=�����{��%�U�����*��i���0�_7č��1L�� V^�W:��5�ƀV]�Ź�E�:�;`�� ���%ofkX-�*nZ1�S���{aj����/mP���ll�̉��9��^��9>��.]Qn�̯
��7\xw�o���L���G	���5�Ƭ\���r%��@��<)r"Oz�E)