----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    10:31:34 08/02/2012 
-- Design Name: 
-- Module Name:    CPU_DDR_FIFO_tl - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity CPU_DDR_FIFO_tl is
    Port ( clk_i : in  STD_LOGIC;
           rst_i : in  STD_LOGIC);
end CPU_DDR_FIFO_tl;

architecture Behavioral of CPU_DDR_FIFO_tl is

begin


end Behavioral;

