XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���q��"}�m���!��g�  Ӝ��$�_�[��-6�N���@UL�7Q�%�k�Qw>�!�vo�&0�=�Y�m��4k��a�]���?��E<�	�R��-�4�tie�~���MJ2'	HZ�9����Z��5;�9��[C����p:l�0�C$i;��/�ޔ��i���.�^�e<T��C���EN�:�;�yiuj�{:��,����^���N-7|���z�HKcr*1Wj���1�]�Ts����C�,n���_�}O�kc�h�@2��=���v�T5���eηV}��%Ӟ &�XwxG��j�sʦTa���Nk�W <[�J<8�����5�d���0{�]�Dy��mB^*V�R��C �$8�rjkil��=���k��@�ߛ'��;շ���&�}���|c�8��B?)C�5!E{MѨ̜��vs�4+�b��p.k<+���,W3��#n���L�!��	�I`�&%��m|�3�a1oCB���o��X�{ߙ
���ʬo]13v��?8��Aj������> ^�n\u�t�9��Rxh/�W�S�h��y-9���Y�Xt�������������i���yd ��(J�6}�������'yW&�y.j���4���֢��?T4f�T!=$R�]�$ڬV�h�a��9�=��m̈́R0�y�C
1R�R�U��~D�xHm܄���	��o����(����3w��<����@���^��$�K��1�8>�g��'��^�ZXlxVHYEB     f7d     6b0uvMp[���[��%-��4��gq�B��G���UaA���JA��e۶8���U��b%epMڵ���i�`��E��"bӔ��;2�O��ʮjr�a���R*M����.�]����!;J�0k\ aҕ��U���;anϖ�ƺ�[)ɀ!]�
����}9��>(ܪ�hUø��L�B�YtŔY[�`�,����=	G�%�R�6A���V�u.�t����3�� l��ǩrF���|��g���<	��VE�����c��C���bz3iX�>��i�"��-���~�;�uI��z��0���9!��!jP�������q7�<��[a�3����\�޻���]�����d{��������?���L�5�Q`��X㚹�`�Rt�܃�ja�����O��Ɯ6�a�留�����l'_%�n�|��cZ���]����������6�;����c;���ŊqiC�9V�]aa��2ȴ_xB��tf�*RK�Q�T�9�'j��G<��D�� �`�!#3S�L=��d�@k��!w�eA^m�3��ڮ(���7��9P�3�h;�S���������!�pǚS��B�$�W�B�?�yUn!O��=΀�ړ�!t�;(��8�"�oO�g��D�+L7�_���aL�YR�C���h�� �0Mb�ֵ.�����8zM�9K�i�gVC���~¹B�n�sdF:tW���fc�y-����}���&'F撀b�'8���e�p���|Rr�C�ڃ��I׌В������S�C�'�%z:i�T	�ǜ��#��ZL�v�T��\������]���o��%��zD��녕��C��H����8թ�K���}�i�t��{p|?W݌��,h���FL.䥼>lIS�z6W��Z���:k�ҳ ���]|eM���<��U������[ɡ1�W��Id��C����~�i>	@K�g��j��|5�!��#И��X����G|��F}�+�:	-���$���dVi�7�^\�c�����C=��u�9q{w�E )yhVr�'#*���}�ip"��~�)���A$��=���GX�JX�w���<q�+��LrNA���ә��y�Ȃ�9��x��h����Q~ mI�O���o���y���	}#։K-sy�n�^	X�����̰jhZʆ��?�8"1{�3/NV+�ˠI�i�;�շ� �ob�ס�T�$�4�y�gHÚ�zH�j0��ϓ�(!b[m"Ň"N��֨��*�C\o�]�Yʯ� X6�ur�E��W ̠��	l�ݢ�j7}�/��E��:"�ɿg3��حZnZdu�4񺈮�`!>fݝζ�m[���q�8���a���F8�`��@��d�q�#/;��Hzb)K5 ��o����au��fS��j��s�_��,���+�x�fV�d��c����i}}H��%Q��
�9��"kج�İ9�>-G��~>�.�9�K�M�v��K ��M��A~��t�K˘�� �����Y�L���)�pZa��S�L�'��ӰI�5��w!����p�v���~f"J�M@%[*H�ZtU����}���:BIB��b%c��T߂uI������
�ã`�3��׋�g��_��7��?��7�n�!�q�ȄA�0�cًTY@�T��