XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���E����v�HQ�G-G�}�XJlUes/@�Ŵn��K�+��@7zr+j�gّ�� {KB�U�E@n�HV�$tqRP3nɲ)�#/��r��SԿ�c+�6뫏�i8�q�(�wѕ�S�V�qLOc.��>�G��*�&fP�Tv�1�h��mnJ3��_�����S���7����'.��x��L�����}wQ�o��	u?�藂2���R��$7,1��d��4h�����qT��TLw�KLfk��^*�:�I<v�CU�/9�/~z��MP�$��p�b�b;VA�+R8��Y�v_� p��T��:<H/~
��^ �l:d�p�}㐽_�g�{�\J��H�3�WK�u}=�����������,>��K� Nƺ,���f`�yIEϹ�5�����!�� �ה] 1��ڀ�L����[�DOvG�p����"���H�U-:���oR��bq�jĈ(2�F�v!+�ڡ<�T� �^$��o��a�߈��MH��~:� Q�3��,#q;����?i���Gaa��H��z6��)V<�7�3چY��� v.�%W���Ȣ��ێޞ8
���%����/��������X��1�ڗ���#�^Mw�u����]�_Y�����e@ʃ3dS���4�p�o��H~�F����or=l���.�Nܼ�b_���L����z�b��z1���l��`��V3����F��{HC8`��/�3�C.`(	12�o��ϻ�2���m�y'ZȻ�aXlxVHYEB    7187    10d0���\��s��!*!8�ղ=��g�iBLB&1�h\�܋#��ۦ��#�����3�ߠ�eo��W��u�7XIw�as_�OM��2��B�x���UnCs@.ݜ�k�V�m���܄��E����T_��?�}��ϙ�������+�DcC�����@c��<��k���5$\4�m^vd�7f]g�b��k���t��
�Do{�����_7N�`�EF�O����xv��{)�r���D�"� ��3h.�N? �%Z�^
ae��������z��2�.�H?a�*KI��*_�-�ˡ�'3E����E�����������Н\"W�Q�w��w�:`j �h�P�7�L
�}4�G�y�l�-jފ:�س�P�&!�:�7���e�'3H�{�`a傥��VCW4',��ެ�ކ��o�Bg���j�����|傤��My�dɗ�T����9�ä�x^��X����/Y��ˋՀ�R�ݼ���rGƩ�ߔ��	/��}�"o��o%�o݆��b��oA���ɞs�EB|x29����e'i��*��iD�L�}x��������(�6�؏������2��L�m1�'�L؉��2 ^�� �Y���l���?u�7�FT�����2��]�N�0�Ä���8�6N�%4v4\+�M�ݑj��+٧{;�b[�<�(p<�}�����;�a���K�"]g(SI/��?�R̳n�w3q� �KI��٥Tl��ew��q XՄ֜aF���z��zk�c5�����:R\M�wR� ]@;I�r����%����>��R�b��\#�e�߭�8�Uo�ma|k�P��׋���e}@Ÿpho,4� W�X�OE�e_����	l��+��cG�'�tau	�7��sa�𴙽_����>	y�
�b��W�8;�VÈ�q�b28��{37��2���ZL�Vi�:�_�q9H�c��/n��9̄�[ �C�D��ˊb���l��u��>�"�Zc[�-Qâٲ���ʇ�j˂W���{Ӂuz���Ϩ��G>�߆��c�vbL}j�&�y��,��^&�Oǎ���� h��vxNQ�sr)��Б܆�����0ɂ�pi�1�8�V�5\�ԑY-R�`�����\�	[�vevn�c���(��K�4����i�-�!a�S랚�G{:��{�tc�2ܞ~Y	A�'�t��@E>���R���Z������S��CQ�v��ٸ��?JH�X��X��.�C�2R�]N����{!A୍�EWFށ����\�Q|G�&�]�/�(�?�y���@��ø5���A �	�a��ΚWp��f��׽��C���4����6bf�$g�k1!��tl�X{n�Z���CwM��̗���� ��˰d�E(��K��^M9����\5�2z��'��������{w�k|g�o�oe��EdR�?���/f{}ӏk9�6ժ٤,s��'a�r�H��ט���4�c��`��y%��M�u¬\��q�����&��M&i?#��'ʰ��cT��.���)UWL!�p0�� ?p���2�8T�%� 9�<��C���ߏ�Q�@�m�^	�q����4���'�?Q(Da�~3����ݕ��h�Ǎ�(u��Ԓ�טj�����ӭ2r"[Zn�D�y:�|�AM̦����e�1�9z�`!�*3��8!*<����8S&���)*�ۛ��(�a+���|��*� 8Rp��*$�d�e�<6�?���9P�)CT�V��9�,iU�K�'��P)����[
�����\ߜ��'�8�LޘQ�4b����GJ�����-�#�����
���(�so!�A7��)���f����wyz�y�*6���+�3RdևT�i�O�!�"�W���Z|�S�i� A�4���8s��:ɓ����w���&l��į�Ec#E`�4|��#�x����%�ɂ�WF�BRDë�xŵ�?�v%%�
o���nJ�s�|�h(��J�Φ���Vy��"��k%j�6�K�HXE��2�$�<Mu�:I��&��|xc�V���O���Sz�z�:��4��F�C�[h�&��[�A����?!q�tp"��1�Q=OC�2��fM�x`Gz�e���[�n�lU,X��CC�x9ϦJxð�|!��X���^� ;�1���<��!+�F,|��=C��q�_<�>��k%]+�P�r��M�Q����^�D��y�������У��x-�bǕ\<o�8������|���8�����c�o���wrflE�ߑQ���1�D��ݡ]X�ep�c�nO��
�tHT�[�dǌ��*3E=�`g]ݡ��q��쫨���\�����H�RR.L ��������z��u�PBQ\_Ɏ�����a�y�}s'����}��]� ��jg8��p�R��fL9��kS�-R�) o)
���8�}W�8=��qӻ�h�;=��h�s��w�cu�j��6��q�\���,l!m ڎkk�&�	�!�z�&�����g�2H���u%��FR�X>�¾�]J�#�_@�G���q��:u���~D"@�p��'�c����qg��G�
ˈ���EX^x�ߺ8jE~��:�NL%�j���H�3�o��xb���2��&S��Ho���7̛I��$˯��5�Y������Hw븘��?Q�o�Ԓ��D	D��=�ˑ����f���gYK�\&lO��)6��9|����B��Y܀�0hqԭ��8�d�Wԧ
$�n�F�ʸ?� �0�t�;򜕢˫��9`������xG�U?��@�s(k+�e����D����w?SM):�(���ۼ�$����>� c��:�n��n��t"��
Er[��?~����-�ڞn%h���)�8 ���'�V�C�RNb��2����:��%>��u�y@���M4���p=A����:R!8�7���%�O;��Y��8�A�*��kk�&�KU��`������?|��E&LX���72���~������Q˸�I9�R���;-���;�JU���:nP�G6��,�7����
�8�V�Κ)(]�L��-h��RE���|�����"�dg����+Pm���B&pT�r3JW��.5��Ў����9t5D+�ԟy�\���4�蒣����f
��^t�X���O5 W�g�32!^$(��|�%�N)X�H��lvY�������f�4Ե�g��4�q]t q��=/����Y؟#]B�?|~2s����q5��ز:��l�tbjZؙi$���jU0��hv�x�?��>XA#�Z���Z�!�����h,���;���Z:'���[�Mfk����9��"=�:��	1ZhQ��Ҟ�j��C��G�G�d8����HQ��#����Uc[vɼܩGN�V! w�qec�W#j�D4�� ���H38���Zė0�/�^�,��Y�oǩH����Bk�U7Q��
��b�)�U���"2�T�A���e(�w(P�w_�U�1�j+�^PUJO�RX^�l۸9dG=lWxOj�O�S{ڬʼ'K�?|u~hRT�\� ����\�T�j�!�n�}8;/�Rv�$�.�o[jչ�j#+;�U�/��RZ�s�����������gk�1�����gk�|ቜ����"���4�r؟w��'](݅�~*�����v w��2�J�=

��%nI]�zu��`��|���a8�����ESog�N�U���{�c�����6��/�<��GaH;oq�w4�ۢ� W�6��`��0�^r�O�O��w�e �) :������� ����.�+�>�&�^��{2b���3*Oo9�xK�*~�ȵ�bx��͚�5����+�7�ظ$� MUR04ew{�1ɠڠ��%GL9v�wߙQ,����od>w��~�"&Jw�$�
�z��eU���
:ӝ�T���H*%�����ܡ������oW/3����)甆���p�q茊N�n*���[�ʾ ���[6� &G�Z���w��b��'�������uD-V^ȘǠ>m��yb�^�����v4������Um��U�o1:�Q��P�����x���
�n��<YJ^��aYVLO��<RF��;]�EFY���,N�qW_�(�����
��I!b�,+�(��iYt�;�"�����������n_ɷ���jl�Bo�Sp|6	]���7D�Fdh�%�+��}|r(�bp��B�(�	�e1o˞M&����	��*������� �e�.����7J;Y�d���J����y�z{-!*�M���i���#�