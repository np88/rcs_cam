XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���N��1�7jh�Xt�H����8�n;;{-�z���A[lRF5AyeM+�H3Y��E�R$Vf���;#�o0�_h�e(��o-~���h�Op
�KG��x� �Z1Zyj��J%�3�qEL%�H.5���AE[t� ���*'.�Vf��F� �����b/b~����@׋��6L��5��lD`ꅳ�[�r���~I�� �c�Ѳxs���%Є5���i-�)���ͪ���$��}��^����AU�2�;&~�9$A͔`��e�  v��`0	�� �n3fo��>�{r���pO1s8��'����z+����]*�k��Q��]����'��:
v%ܒ�����8�&����ͺ�:�i����vX��;*�'��P�J��o���Ei����������>���tg�I��$�+��r��yۈ؟��2�"ʀ~��4ȁN��[k�j_��S夛$�����-2���S�+e-v�is��n�(%O�
���L��E�}�}�����@��V��ԩ'0W��gC3�;�(�+x�������m��$g�T�`#2��?��i�'��`A�}&�~�����J�6�_I_`�'�G  (�N�-�S���ŉHn��d�e!;~��mP��!��l� ��.$"g~�K�1���{熛/��<ܭ=�G"��]
�q�� :t�<6I���>�%�OÏؑ��[�������z9�����" J�
q��ݳA� 4T|}�HQB�"��k4XlxVHYEB    5b76    12f0�DO��}���ߣhD�kQ�=5�7�`�c����nHuj�[_�E|J| �{um�ll�N���L�A�kHʽ!idwS�����!�%�o�)".ց��:���=���hnf�B��� ��`�}[�Q@�& ^�'g�1R�����N{Pꩲ��0?���^�:��=�5�ԛ;i�q�3��� h��!SDS�1�O����d�	�5Q�N�! ��[��r�۸�)ˍgo��$��A�cʨK�ulok�}��e�����[�P��!��-� ��7��\�:�nC��u`Ō�it� �+�IAUG��qc�P�B#�ܩ����B���"����Ѥ�:?&WŒ�H�xI?��<M����3�)�ց5C�GS�]�޾0�
�\�����i�N�̠�GtNhu�\�%/��"�B�,��}l !!c��耉�gE�Ƚ[Y���a� R��$�0��p<�d2@8�J���Y�<q&wSvJy�+���P�ݜVFS$K[����2���&��5)�&Νem>;	��Ҙn��kn0ۛA���>U]��.�T���U�<l����hx��l�/���
���N*������b���G#ݛ�R��%�`@N�{7h�^�j�m�4ެ�t�8�,zR�Kk=���V�����wZ�]��p<6�1m�}P.�*MU�zY�e-���k�XD��bK
c�%
����"c R\�+f���?6��)<���|>r����7/:L4�ǔ}V88 ��/�z�j�!#�_��}'����&m+��$q�JJ_��'�&0��v���­��K�rv��p�R|����%��**�g�f���3�,����j�d��:6t{��f��i 
B����.nF�Kb��0�@�AM��;���56���C�U�v��b�R����.�
f��p��ح��Q�d1��f�|�+� �|�z���O��)���S|u�vD�:Y[�v��t���&�z5��į?�
yoEU{Xv%/�~ّ{u�7a��H%2>[j��ܐ��N�Yj
.�v��D�w]�˷��s�-���Ni�~V��!�Sv�ĭy��sa�6�P��P�H�2�#��T��W(j:�E��K�|ƹ��C��:*����,��O�1�-���NM-��z��}u��^�ئ�ڥψ'sg"� .�����(>uŽlE9(�A�Y����`,l&G=ݒ��>fo���k�\�Y�O6�q��8>�Ǔgj����|��'F���!�9��^]�\@~����6�'pNx(����Csyc����j\��%��N�:����Ui��XW'��C(�=[J�\�9���ff��㔰ԡ\̍�ɥOE.L�+�����,v\)e�zF�EI�(� V����[����Ġ����)KH�~�x�"(ŋA]�ٗ�P̕�����Z�~Њ��tJǪ'(�kd�SY�(j$6����І�}_+&h7��fL\��&u�"�����D�)���垏eݺ9d�g���/�-9ED҆�"F� $x>���ZBr�ѓ��m���X�T�+4�y�-�(�d~<�*Q���'����e���qe1�d3�~0����m�b�d���Ԏz7G��7� '-b�d��<���	�R�gB5�f�?��9$��@rG�<���n4	�h�2�juW5�8��H� Fb�Vm�PA�v'��\P_����XV<mt���'����( ���M�v��J���o���Ɵ��F�d߶�̎��ٷc�9�JW��({֖C��^�����|�1k�lUX��-s��{ߺ`;��]q��(�8�؟?������8b�>���NmKnCY��3��P4ZǠ��;YLv4H�0!	^��r���a����G3����JH�Xw���+a)�#\TC�I9Y3"���_cX6�L���*"Y��Jt����^k�Q+�!mM�/����f.� ݟl����q�á9�K���~�~\�B�y<���Y([�����m.����6W��������J�x��u�5��m�#�h��G(�"ɼS���
�
��O�7��0j������q�5�ӛ���r��;N��θ>�^[�y0�������}%7��5�WJ��)P��^X�_��B)����4�ͫ������bj�3<�%�beAqSA��H]������&K���}�����|�u����/B��|C�>�~��V/�ſٌ��z�s�u p��l�7Γ���M���56I�o�BI��`1sv�1H{r#/)��-�qj���z�#^?=.-^�a�u^�A /\�&�+)�Rn�䓖n��V��zf��G�U�K�u��.����rui�C�?�͟��+̀��3��7^��N(����+�kn�ń��i����z� 0�<��O����A$!o��{�ۡ�!�KA ������Ӱ�yNJX��e�Sb3J@R~�L��|�)P�F�}m��}��w^�jc8p Jc���P$'8(p�P����V0#\��`�a�D���6�G��y���T/����S�#��ܻ����#��:BɍfIN�Mj	���]p�����v�tD��xa (��J�B9)����>;F�����K��eo˴�v'���{�n����n5�0�$D��=(��9�P�B�}����/	֞�I8�?�V�ٙ�}O~͑�'w�'[3X�z$82���ҫĢ=��PJ�=�� �̺�=��U	ͻP� i�!�ߗ������?X�R�OIh�s�]�L�3K��f́i!۳J	hO�q%�פk	0o����V��.K���u����h�J�T�2n�n�F��#S��I�x&��wk���lȭ[�`���?���E,��g^"�q��`At�b�e%�o����T(�&�߭�&P:"������-D��]��j�of .�1�ФO�B,ʯ�\}��TK��vC��pnEJ���2)j̃]z�A��1E�Ӆ�H��${���s�_D�]��Xu@)�%r�M����c��#���)�D�N]�PJ�1���
��8>^�-��y��:�?�cT�`kmoN�d �Pa��S�N._��A�V��N�Hw�0h>R��qmF|E��2p��36��Op��{���is�hZb�\ �pl; ��7��ɉ}0i&�BŶ�\N�qXl����#���Tp����NS�*��$=�����fN�ڐ�7	��u���.�{��P4"/|t~d�_���e����;	;�"�C�xlI�e��A�9>�uo�&M�)CQ�Ybn�sÑ�DWqN<��@J���`7�c;����8��?�Ň�,�d��6��qBܜS"ݼ�P�2�e�?�
�P��*N����wH8�JF`幈�6�!��۱G<�Ó9Y�,��g�5#�Q8�`�􆈕tp�6̃�|��h��{8x(�a�C"p��W��t�>�øGz��M��w;/*��5�5#�f4��ƻ+˴-�W��B�<�B|/=
D�b��egH#jG����񡹹7M�@����A��q��!��Ϯ�+v`����k4��[-�Pn�}+"O����.H��ت�Q�Δ�H�$8!Ys�ɡSO�?���6���8s�v6L�K�`�j��-\)������h\��C�HDO+COqG�˥��B�U��&�p<�~;���m�;�3"�qL%�N\wޘR��; $�u-Q���-�V^NU�3Ș��A-�3H�0��{>��Z���%�n�\��F�"仌�!��V�3�!�Á�E�u�:�FX2��&@L���>o_`��oyToJM�r�yď���
�?*T���yB���+�~i�F	�>�`�(Z�/�����G�h�c,���mf"'��0��,�#����\�P�g�Q��@��D� ���$�&�05��j��\��C�`�NgF�f����J����a�1DjC�h�G����&\,t�2�/Nm��Bfz�D{;q�;�MsT��snmf=�H��^
�a�%%��W-�¿9�r�y�Wt{POyP�#A;�Z��c!#������?b��v (OҾ�)���X�8%��dT[!�G�h2�K!��ch�������ƣ}���l�Qe��_�̛.6�)��!�����x� �c�z>I�W��c.���!7�o���p�G�-���0�d�*�q�����Fv,һ�՗%tdU��5=�;Em.?f�eŇ�R��C�죃1��x<�x@���iM�q����&�칸kR���)H�uP}}�U�P�.P�M�J��'��Ԁ�Y���A�Bh�=�.W���P�R��^ǝ��A� .x���f��([I��z�R�L|���\Zc��>w��D�u,�s�`iO5>�1�l�C�:(B`�3���l����'�!��t��-�ex3EZA��!G/.�����
!�}B�Ze�����i���.z�M�f>���B��'�uLͽ9�\sP�<�N	��FpI��b콛\	-;�lE��!��+�n��w��+�/�G��;��WB�5,Ţf7ӕL��kb�u���L"�E_JQ�:���6���" ��ң@�6�%���|�A=}���b�$�Ě�5�$ aR��2�x��O7���`I"��00��x~����D\'��ץ�Af<�^�]o��n��M��Q?9M�p���F���ӿ?�3��{ᵫ~��a��{%ͧÐkʎ�w/�j��" ��~��V�xx��#-�{�Q�K1!�yL��j�=�$�r~�vǊV~�H{���W7<��隘��o�2ۑ�qi�Cx��n��^f�})��Vf�������RF ��XnF�طSJ�&�%�ꫂ