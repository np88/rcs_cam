LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY Microblaze IS
PORT (
	fpga_0_clk_1_sys_clk_pin : IN STD_LOGIC;
	fpga_0_rst_1_sys_rst_pin : IN STD_LOGIC
	);
END Microblaze;

ARCHITECTURE STRUCTURE OF Microblaze IS

BEGIN
END ARCHITECTURE STRUCTURE;
