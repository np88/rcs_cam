XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��8�$,�W}~����@))���@O59l;�~��
�I8ؽu����-_�,��u�_����1%��h�B�=_�9��7�GԊ�NX�����5���S�~��c��I��}��Q��S9���{��P�	!t� ��f�Ynh��;����R��ܺ��|�FϪ�԰͠Ӥ�{(:9Ȥ'���c��x�K���(��(�[<��HA�B�E�K�������Kc�\�2�/�����Bt�L�|<�����͗K��%��E�/����z����2���@�bE�daY�l	�[#�Ŋ�g��a0ͱ�\E����2r��;�e�<5�In�����	�<�He��-��̼] ��󸽂1�`S��g%�"����k,�re�i;���JQ�y���5m ���>�(3f=bcGӁ��N�Y�0�3�T��}�O�w��v�BZ�W做��Ó�@�aA���t;����*��G�0���=)J�z�{�2efa_����HЂ����~���jT >`�3]��qqUd?n�2�S@2V�	/'k�L��2T� m�o���|0��Q8P�S�.4Q��_P`�~�iE�y��gx�PĥRM�=d��]_�\�1�U�\���R{��R��-�$'s5Z�$��O��;�� �n��n�Ew ��{,#���°�R�T�+��=�3�����t�xv�}�Έ�;�����(��mȪ'���Za�ago�imQ(Bqg0c���ܞ���{XlxVHYEB    9193    1ed0��ĥ�Þ����I%��;��c(�~ �������>�JǢ7O���z>��[q~3����%�e�!kp�<G�W]�tdn��)p�xbr����7m�ʘK֭��W3��<v�Vg��:W�ET���]Zs/��-ҏ!	���J�(���A_1[�*�	l�S�Kܞ!��A��ԻY~�\Z(�=�c9[8:kN�y��(Fz��qW0�/J� Mt��o4Q�z�N'���m't�v1�W�c�Ja�ĝ��b�����ߦ�jxXR�t~�֬:�fw���6Z�0�.��c�ZTY�Ra��.����A3;��Y��r��u����zY��0����J�����`�θ�&��n�f�LB�K��C���%�. ��1?T�����v\�_�A�S"��!ʻv7d.��A����8|w��x`�q�m�m~�|}�g��W\�)~SfR�o
�EGө�r��X�c[�bWK����U��ҥ�6 �d��4�\�o�4�	P����=/��P�T��[*�^6s�8e��}E{��Z�im�?>�"�s��k5b�;1l�5�f�YIˎ�_?�#Զ�p���6֕�3��?��N���L!I�yy��X[�~)��ZP�u"�i;�o�0X�5X9n�\9����WY
��TL��4a�C��YLo=���o�������=�6|'@��dW��>W��es�3H�`	W0���W���I�=>a���R�6�v��B�4�z}Ϩ�T��u�������5L��g_:�����zL�m��N~ȁ4�d�����`�R��'�j������R�Z�0�=��4਎�p)�����R�(���@5�2p����+�nё�%�b�ˊP�V�4�)Ϯm
��hm4����G<�O�2���#>�s��u�U+O/�-$�w���m�M3=�2�3ĚU�O#��Y��)wpk��Bb��`���ͮ�[@>�T'�R�%(��pQ�"��)�5��Vj��j[��,����j�rq��q�Bۧ�}���#�xJq����y��]]_�jz�^��5O����9�v��Q0t _��_αȞ�A۴7R��Bh��oxe<�q0YC����_���h����s�$�}�ب��T�`X'�V�&���/O����P^��҉J���6c�=�����I��jͦt�ϼ��2���Ck����q�����-8�I��8ŭ��VRe��d�`	��-2ⷙqR��7!��&;��
�O����gMf�c�֘g�Ǽ�Yz$��#<:����4��!�ƒ�#x��6�u�+O�-�x%�њ��s�Δ��U�/� ��54g��z�K��[�������J�������3����}pK�bU��kI �e�Q�5�;^������/�KoO�پ��9!��|(�yb��`=��f�k$����w1���o<��Q�F|53'�X>[��f�d�Y�
/�8�g����z�і,AY��\\]�Z|ȼ+�^v "�$�;�h�BPjYR&'	ܦ%en$�ω~\Ԏ��sL݄n�iL�?������Ӟ�;�dǶ+ɔ)�u�!��SSҒ	�/B�U췆��)/�^�x �G`�\��fl�ҭ����7�y�d�i@����`|�Y�����I.Qj��^X�����oYj���9�KQ�FS�%
c�D�$�7
+b�LI�4��1sK�.[N������+Z�����竑<���qe�k��u:2�Ճ�1����j��SÐw��ܣ�ch���(Sl�S&�m��Z�:'�������h�H�)l���Y�\�R��;
V�nЉx����q��<h�%D�X����?��Q�7�\t�c���B"Hĥ�C�%ª�ۊ��A@�ݐzo�I�0�˝��Z|�l#)���\[WH�t��x���1"je�N ��g �,Җ�ѥ٨�|���v��n���/+�&U|�^,��%t&����F�E����\q3}7��2AS�A>|�z��$��<}��=�Mn&�Rl8rET�am�1/C��"�+�l�!t%���O:���Vw+U�oۅ��"�{1�(�_��F	�^Xsl=�
qKh����k����LQk2,J�t9�s�
X2u���(�>6ʛ�k.�9gҺ�.d�s�~�0��6���@U�e���x� ^ �K^���F��A���+��E�	�n0�ke���RB�����B�=��aj�!Y�&9��dj�l6��<� [���?�<#�\��4�W�11b�xPo��e+����\�#(��j7fÛr�c�ZlS�D�b�G䈵6*�'���z��<�t�UZ�E�&����д��/�nΉ�u"07>֑�q����C-�
, �*��;$�A&������9����������Um������յ��iP�m�U0�ܣ����;`rt��'Y����G��k#���������'ta���gU�/�}\x�����#n�(�ѥ���b�Qp�������p�q�@�q m!	<�%Œ='Z�����4���Ĺ�|�L�T�7�Mo6��u�$�sG>���4W�='N�uM�\6�����������Pi]\�����k�)x��k��	��2�w����h��J��Q����x0��g������mVKqk?�-���P��ZZRuĔa�����f7�	�ҥ��q6ǚ��-~�,��}|���z,m#̛�~�AM�:�[B�b/l�sN��� �Ƭ�s��s1��u��*#���0L�����U(�@�p���`縪~�:�H_UT�>����e^�E�7)�u?u^ћ�� ���:� ����S��vQ��[n�!N��N�}�ϵ�m��k�mB�r`j�Tu)8��:�g�D���m��1��<v�X�[L���+�6Tc�/r�d<������o"Ü���3Ԛ4�m���E(-W;����-�^���S�?�<��:��U)�#x�'�y�Ĵ��5���q��<7��x��k+m�{�VM�%*5�0u�y�hC8��Ҳ��cI�������?FS��#Cr��E����%�I9O�G�tσ\ `D�җa��:8��´ m�_G�Y��n�T�0�jn�`ߔO;�M:2�\�T�}.d�̩G��yp��і�Cͳ�ટK�l#JH�`��Ms��Xʚ$aK{ϱ��jT�IQu|��F����(v�`�����O���LnE�!�C�14B^�z��)AD=j�nAZ;��O�=��E@�O �m�<�{�Z�s����S�x��rP��0�IjO���|�0MC�(F��]��zbg2�[�kq9��KU��iKD��
g��M )9?A���S8���S��i��G�-��>�B�++�.ͬ�1��*O�4��� &�-ߝ#��c��{;��y��߹z ���/�8��e�4��*0�J3t��w��U�]�g�15��!�Җ4z��gތ��I�_w���{�c��z�~ֿx�/�S�_�c桬���!���e�ȶJ��5�!H�e�Y�������E=:�A�	������=�]�ե!���� ����^25l�E�|�S>c������K��,�k�X���ك"B�J��`��mW�S��`F���q�_s	�A�l o �0ty��Qt$Eo�bpO�i��l�Q9K��@��a(1�FڻY�U%|��P��&���x�p#,}�z����ﻏt��f����a�ӓ 5O�s�Kg���E׋�ж��|c�̓��̕2t�}VN��'6Kl��k�JJ���=���_�J���֧D���*�?�_����V�V8�	^-j��2	kF.�'����	Nb��7lJP�Vc�.J��Pw*��	�E����}T{�[4+�P�
#�����5���{#F�_�C�-_DM=���L߆�Mb>�׮0_��&�`yZ~�v�s��m�5U��o玡Q|���3�I3�MU�,���C�QR���d-�>fI �'��@���?UEZ����N�[�M����f�S#':�hF~]��?M�����<�Eq�bP�ha'UL=�wN`;�>�$����N��B�4�N�r�H����"��J�(�h�[�l�r����p�a_�)\�g�^MҫB/ʟ�CE��aqY���L�i��` �>����vD8]��z��M
G&�W�?����ު*���9����d��<�̐6�i��Ji!Ό���K�<a�2�U'dŎ�i�V�V��׳$xeg�Xkf�<ftS�c�TɷMY5AH�����M��)Y����3�Gl�1�qt�,�yz$�L�c�@�č�s�:}��pȝ~p���L�����؛����
�]/Q?;=|�S��ޥo��J��<�c �(T��&�Q`�Tug���u��@����2�jF0T�t���Mscw��9\u�1.R�;�j�&�R����YA{�..�7��Ȑ���p���ow�%�GM�đ��b�f�_Ufh.�
�����Θ����*���)��_�ώO�r`G_�;����`.�a�~~HX�}���҉%i	E�2_��|tڦ�²�,;��Ģ�,�r�(J��t��	��_}f��#>�,�6���@j�>�&����GZ�{q���5̕��n͘��~q�:@3�B5un�Q�a'dQJ�4s��ʆ��V���1(.0|�ok����]d�6�I��i�ŝ�����f��|xxfT�����I2��omH��l�ǲ��F�U�-����/�ԴF��휏v@0��MӦ�+���-�HhrQ�_Pg)���I��:J;�l8
�KƠ�`�vQ�P��$\}�P�^�'��L��~��Nrm����}5����V&�?7$p�m�����1B�u3�p2��ϗ�Ǯ�kĻ3[R�ب�v�ފ��m^�
W�W�$m���6}71�q���_���P�B(�"	eh�*S!�}���a,%,���s��$�ew�R���"Q�y4'��I1��T�?p���L��\����zh��{/|��.5�[�Qm��qՀޖ��ػ��]�u�%�暓�DI�}�_�lj$�^؁WDW[�ZREڞÅ�*a7����9ƴ��*�5g��V`���R��7(n|��Ke�@�Y&Σ�5�a2&]��7P��}
1�qhA���]yp�\�ˣJ�:�*Ŵ���W�|��F$���n\��/� �JM(��s�(ڳ��:Hy����ߩ�Z*i5�|{��Q�4ڣ��aH�mTI�Ql�#@n����d%`��Y�I�%��%E�@����w��0zd� �����Htb���"V&�ud�2��.���A��l�4�\��P<	@��x8�X��7l����
\c�	�Cx�u1������ьm��N��r[K��1�hN`�u}@����7ݠ�����n����qխG��U��F�&1���mڝ(�[I��hZ�����%��E�8�q$<ۨ�nWAǻ�Q4�:5�g�Y+� ЖTs�r�$q�d�NP=���.K��M��mՔ�-|D�T4%	�peV�_�Y��I��ToJA�i2�����2��W�[	�vg^;��r���.�g>��ݛ}[z˪��q�)N�G��٢�1��ة=k�������^	;�	��o�ahsf���~"M,��M�BG�)��q�7'�X>�n����	�M�TL�݅�3�#��5���8y�Ū�Y���˄&�ߩ��g��~�����v
�ل;|9��FB�[�5��d�Zl�K��=g��5؞I�z�wMm�&�D��t���{��@	��k�׮���Z�-BF��ՌM�'��]��ٖƶ��-<����p�\z��
�.9�q��7�Lhs�N�߀)��MDĝ
��ً+O��ο�af�l-� K-��^T�Z<����^~��8���ةh �<�8�Tb�� w���p�m!�}:����k��3�r��h�QV��g\rћ�tu8o3s��4 ��ReG��;�����˿t�(#@v�:��t|\j��U� �N	��S�$���F�����
qJ�ܠ�r�M�LOٽ6�Y�r�G˹�T�s���3�՟�����!c,�J/��D�U���R�L��p>vi:��1;o���b���$Y����d���*��ܦ���t>�I�N������^���:.��?K(4C���s����h��h<��gU~S+�S�Q���~Tw�d�r8���xuM���.�n��$�X)� �XZ�����dQ� +��P�O�ڤY��;2˅�/�3p�Wϭ����*Q��?�]N$=�]���s���xO�Y��ZR,�/�L��.��-$��z{��I҇��"�/����ޕ�e�T:5;��1���u!f�܅���i�w��J�G%=V-�m��;p�b9�P T�1��s���r�чЬ��c4��y�F�W�����H_ĸs�=`T� ���
�(�����B�8�����7�k���:lM ��V���!
��)��3&���si�b��ß�	���C����^k��'8WQ_o�ZTm�W�I�{�{>��+'��T�̓���R�Y�CC}5t�9=Yf�Tb9�,��d�o��py��[��sX�� �5�@zXAq����gǦ�c���G�g�)��'��z@�:�w�rM����(�D���^��C��D��8��ր��XH<G3�(q�ET6�X���+�)9T����I9h���$,�����Sh�~x�[�Z�7yW��i�u\"��E�a��Sy9j�
Y"y�Ӆ�`U�O�CQ�/�y�+��s��3�z�n�e�u�P�0���·�a[��@�$��|�/���5����M��-h�6-L����[��N�ᚇ���'�{��I���..f�d/ �i�dԑy1���Uo�e��Y{�|T�WA'�#�So1)
+*ZR��C}�-S��(J�QL��p�������9�Fh���S��F���U��Vi�v�^���&S���7
��<��7^�lp���usȃdj~�t��|���b����ᩔ2F%H�o�ӫX�놮-u���ȁ'
�����b�ӧ������e��(�2�#�A[2)�l��,x�	�}�$V�[���{�/Ę���+�
��U�a����3�/P��cvra��]�Af�'������RD�	�hu����F�`o� K�/�w*
��E��A�l.]@�I�Լd����	�{P�irw��=����x`��Z�M�0q>�Z"������O��!ș�K���6�~(�ϸ�MS�D4��C}b
�5�9�vm�q �L�AZ��ݎ�Ln|Ȃ���U8�e6��,���3�D��a��We�\�݈�THJ���B�cm��\���]��.~��� f��,&{�e�����$I��)D����cק~�8��j+��M'`�UO�,�YX@zr%sА�W���&����g8$w!Uեu�[Q
�V� �v�]$ո�9� 6�)Nv�˪&t�f�#�V�W$�OZ9�V�>^�>[WJ���ffwK�}�gɧށo�������a,�t��?���S��y����癊?���R �w!����hҼ���+�)6�>O^XB��(�[���YJ������C��jE�LC�y)�=|=w.F�d�Ʉ���~[x�6�5��w�mp.�n-v�����:?��ԉ��*)���j��̋	��>��o���L�ܱ���q5�����v��4���؎8�S{�JVcz%a��&#>��M2 E|��Ҫ�@���|��WC�Ջ���A��)\I���