XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���#!�D�WĨ��t��ZKP���,��Z�p�p�m�y�����C��
�.�F[Bu�ě\}AU��_`)�TЧK䆱��5?m,ci� ���em�ޠ�,#���/,�=�H����#ƄQK��E$JJ�K�������]v*j��,�B\e�~C�c���v8!M����G@�����mA�P��g
e�Lh�z�*Iį�g�9PGB�v0M�|�'��'�n�|	�:Ȥ����8S ���9�,�D[��πK�"��$����e�_	ED���W��1���Z'�B�Ӡ���q�X"7G��=]C������U����:]_��K���*a��wˍ��t��^����(�)�����7A�+���K@g�I*8*�,;��^����k�C��V�L{�h�����('}����f��J��g�n�p�v�%�_�Z����;i�R�2c�em\�)H��� ���`�Zt����Q#|�.��O�-s����'�a!��8
W�kT0U��}@/��������9hW�f��؇�P��P[��R�	�i����y×���s�bO)�����K��x�:�!������ә�p���=��?�^0�Q���g���b��p��l
�������:ii�F0�)+��`���,��B��=�@�t��7���eQ�Nr�o*Eq��Ad�Kt�<́y�Jɻ��E��O�K��?#ڄZ�S5b�:KG�&T3�qj�]Ž�X���Q���>u��=RA|�'h����:y
XlxVHYEB    4089     e40����|j�猻������Y�r�"7�,�	���E�5-����nőQw ���eq?����6�'��Ϙ����N��	M G!<��.R��2􍏕�`�Ck���I���tF�H�M�@��0���˞�N!)�'TR��F�9�-�ӛ>����7p�ojdR��6�R(�̝��[Z�?.�������S!Hs�Gk/���0�{m	��R̃�\Y�3�C�?]�v�M�91\�������P��M��޴�@�E-j}E��C
���m cO�ŬW ؜��<O�����z�ZT}�gL�：�&��=��z�e�� �"p�w+I�9@C)���I�;�L���(�"����<6u �&�9����}"����D^ux���y�s�X�ҖNe�)񤇎���v���]�)F��~
x�u>J֞�y=|��g�қ"���[�j5��.�����3|��%�|����i'3^ϖmE_����̓�,!O`L�	]o�5²�.m~�X_R��)��)�?Z�L';@�0-"@i1�F�{22��^��#��s�zy����(Aa�s����ٚx70�j���!��,��)�ѿ�T��ƿQ�<Ⲏ�E�z/��*�C�qԷ������r_{w�6�~���ȹ�W�>����q�~5W����y�LɷZȺ��Na�Y��{q��\�|oQ�M݌��wM���xB��uͿF�xM�]1a�lΦ�ץ���h��Ef�iǤ����N%�L`��F�JI��\��OV�,�ܻ�ז��U�0�x������8�4����ņ�+�n}�9-2K�39��$�z�z�%�Z��5{��>^r��N�q��t�U�z���7*o�W�!�DWA��i�
m2 �����Ă�/�[�`ta�,�]3��Zm�2Ӭ�R@�:D��X��1��C����`ܤ�	
b:*�3��C2h�э�Q���Pe��MQ�v�v\}�5��!_L��u���H�(�[W��M��o��@��%N��U�1g�uꏆD�커�E��j��<�'(Of�j�#�Uu���J�/m�ze����[IR�H�0��������=�|�O�d,���^;���GW-�254�W������N�7V(I�x��`n��������t�Ww7����@�G�� ���]��0�!�e9�S�m���R�KAjA1�T��J{ac�c �
�j�@�2Ȃ��As�Nł߇1͍�L�^�P�6��BL�ZQv��4�/pr�h?���� �8H� \P^��V���o�4�B`��Z���	�S]4��%Q$��7����~�"�'1�U��IDP�ouf���q�e�<?���C�yK�[*� Φ��0�4V:��\;w'i�D�0)�
$#�d$!���%C�h���d�^��mV��͐Ѣ�\�O��E�6ئ
3_�k}�=�.�6B��*1$O`�����4�Ў�8
��"7�k�_�P���Om!�V���:�O�5'��"�*+~x�7i��P�9��8ڍ��8z�B}�Vy��k9��Pظ���k�&�]�7~�;_�c�~P�5����B�z��dX���-�rEܪ~[���*�	%r��q"���!Z�E���y�r\%��%#grL���C�缶��L�����)f�&�s
������Sa��A���q0������ ����l�ѳX�(��JCb�8��t�V��N������E�.�J��zoa�]��>
+9p>S��8�P�@S��c@B�5$���xu��R���d�3%E�����ɑ�=.��E �C��ǏxQ�q��T���2t׃\`2�;jͳ���[����\������I�o��ӯ�$�h_H�'��!e2c�aO�^��{9?�߉�e��K$=���Ѝ;C�|Ε�Y�ٻ��LG �>�0�
�٭��[GB3�?h��u%��Q��BV����9l���$t���e31[���P!@�(F.GG%��C�n6n!�B���s�0�U��3�!l�!}�3Ye����9z����S�G�%�#w��q��G���c/�!����;�w�su�ޏ�Z9~A�$�4��)|�º�iJ
8r1&#Y���B|`�mN.�F���sX�n�IC{
0�^�2���Sٞ!v1l`���C����&�D�V�P(i���k�$��E-�=6���Y����Cb�[��:ug���3	W�RS�g�B����c/�9�9�A��?ܜ!p�X~�K��,MH@��Ow�ʀ3:�2�i�';� +˚�fd04¼��Hx��/s�ql�NY�ZK������)٢�	�U�	Z&�?������	�$쵥\��+NC��?7B�m�����*�B�:����c��?S�T����!���W�T������h�=�=��_.�	��ɘ��Ⱦ��	VLҞm�6>�=F<ͨ+>~b%{kvF70w��I�;�-��1�k�`Y�s��=×�h�Ւ�h�9w�D�]���Z�%�����7I|F�QV��L��(aj*��<�6t㨭*��kEz��y<����l	�;	,K�C<Ty�*%D�غ�3�����B,��dDL���$�æ�ʯ�w�wY;�O2Q���KD��졐�@��Ǘ}�����������^]��A����.~��{��8�z�B�8�P0���5���SJ��ՍvO����>�J-ozPk� Uo~�x��+uh��eHs�ߔ����i@?(������Wys��_MJP���>I�����e��H@/-5�)D�V�U�y=3��,�����ch�ݭX�q��$�2d�G�Smh�kڐ$?c���,Q�ط{"a� ��P��nl��C3)2Λ�#�����`���f�|�ø~�����g
�׼I����bЂO&!�VV|�K�ׁ�pF���]�;����}e�|��w���ѻDƶ:a����[������O1V�A�i-�6F�3�XsS�x<��Kp���a��B��e�P�B�",�$������6,�����#)T/0�,q�����4�ׄ�1�����6%�p�ˤ>�����H;�N���#�0��8��r����N!#��Ƭ<��t�V*̠�	�W�
o*ڃM��/b�ѓ.Z���s!,I��"POO�6��9�%^��*ycŝ=�l�X������ @���"Uj���4&��ou<%~-c��������bU�v�2/�l_y{j;��/,Ү��uj�[��\t�ӄ�L9O�<�oy��d�Ș��<(�k��w���7��Iuv�_�7���i2H�K�F~���d�8�B�8�x,!I��k5������<f��,s7���R���� ����T<s:[��!�@|r>jP�ь�Z���a4m�t[�����@tN1iBW�e^�y��a���>^I��u+�B�υ�o�� �E8�p�h�<M�<Y4��,���!��	�k �~K�;(6S�i{[ C���6��0�q(ۘ�
�Rjj�*�vւ�` ~���U�����������`W�n���!���@+��SӜx��Y2�7�2D���2͓|��U�j�e��