XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���Dj�:y�I�u�f�`��	�.Ogh�Qs��ǻ�S�jޫ�7MP3��O�`�	�� 'r�	��~[?}���m����0:����h�� d$���Ԓ{�QT}R���P+�Q��I¥8��ϛ  ��n��Uݭ���Ty�J�F%�W�i��:���� ���Y�+w��w����G�ҡ�jÈ�Z$��ӈ������yhGlZ|l�P�)�/^/�UÑ�{�������
S���s#-���\��;D$��Z���{u
۲��^eͭ����*�o����Q�w������Rz#���`�Lb�3/P>Y+�l����?�ʱc��o�~�͖�ϋ��y�<t�9G��[�o�=�lҭ���Q��"�_ހ}a9�!��=;�{迂W�����[�d���WU��H��&��Z�˶�Y cF�ϒ[���A�l��w0��q�J88q�������~�fMi�e2Y���RZ�E�QԹ�H�#���s�/��nS�k����Y���"��}�����>�q�o~i�dD�c�*��i!���A��S$c�c�6[d�r�)Z�E��~B�)�q���ԍ�c��x�*�*|�o�zw�6��F��Cd����p�%_�0g��pSEpZ��|�y�2��Л��"�Js����5�M�xqD�f�z�����o�?,�"i����U��o��}30>�y��oք���lM��9Ϝ���n�n��	А�����͞��xQ�Ԗ�|�+�A'40�wyW�XlxVHYEB    63cc    1460�4&�=ݟ3�W���~�R�v>�k��a0q-�#��$���]�~e��%��p�-44�N>�aͭ֬�e��\-�W���W��-y}m:p�,��i�y^��z#:n�ֿ^F���0���v��?~�G��#:{�R�ʍ�tA�zP�[���������1vT^2�xu�Gު?�pc)��	�A����|�;&�6�fQ��#r�b�_}�^Ǟ���-w�?*�8,E�Ժ:��|�x�B3cS��t)T���Y��4�6���/C�QN�
�$b.�J�^k�!8k��[��.�L,��q��1�0�Z��fT�؞��4'���7Ȇ�^�U}6˔'R�B��oӪz@ͧ�K0kN�` Q.P޽I^ ]��	ˬV�V�w�f���s��_�x��_ n7��*j�l=�\W#�bS�D����gl��▆�oC&�y	��l������ѕ&EPo�a���M£20d]d>�Ym^/k��~&�/�@�Y�C�7������\�A�=�~�2B���Z8����t�A�	�M]"��C�jC�Q�H��Nlq�&��V]��� �G��W�ǐGŐ�A�<Rh����9��̏(OTV�,�t{8,� �q7�E��p}�g&�94���uHB��˳{��:1:�`<��;ι�����j��B#o/&���5�?^�Yh�8����� s:L�G;;L�/�y��I�a9��B�2���c֡�#���j<bO]��Uc.�Y���y�\�m��~�y��d�^s�=�:ɣD'�3�9���Le;$�'��(s@�۩O�k|��~Jª�A�sF�l�q�n�Q�d�
�I�G3�9���4����}��֎Ӣ3Fҙ3�4y�9�.�:H�o�5-/�.�"埣?l5R٨RPs��W%O�6y�&���G0y��'����N	&­m������]p���l����/0?WD�)�&��Â�����F�����C�Nh^1흭��4r�s�@��*"�"B�f67��4jfR�Q�Y:���	P�m/D�9�W����G��P�T�j��f�*=���?'�z����=�� ��� �E�lV��x���k�mnt��4? ���|~�ų	P��_�	9£3�ܯ�k�5�����a�zN�Dr��d�# �I��\K�����Zȓ��CP�����׷0��Y̺��|�����+�$����/`=�{�jf�E����+�B��y��.HvUQ���T4�O��jf�����c��L=hy?~��T$�t�|i�t2٪P� l2���w;w�H����$�~|�9n\Y$���:�'�����,��1{l��쿿�Jd�o�p�&�9�K��S�Gm�+o41� N��^ �b�z[�u��U��G����E�00Bs"�9�U�dE�1�<�g�W�8�6���b��#UeQ�.�[��*X]���cʿ�9�'j}��v�[,ր��pF6n9�ۯ�rF���VI[#r��ŵ����H�{ �U�T��Ċ���NgN��uL�D��EN����3Na���;b�C�D~|�:{���"7�eƊ���z�z�������ލ�'��V;�_��kF����_�4ߧ�b9)T;��R�#ứ�Ј-�夫�����y1O��_D� F�pܥ�E�:2���q���?�Q�P��H�xE�N0���C|=�p�F^���!4G����@��E�2�q��]��e�6_�Y�R�˝��[�hݦ��h��x���}�T� ��`#l���6�b�ic냫��y���1��潜`�V���w>O�s��đ}q��8��!���P������GR=s��sVOӤ��
k�JvXr[�Vl���]�\�H^O��I(�?�T�-�%�]�!�Z4{�FK�mG���~��޽u�l�K���~�k����C68��'�V/����S
Wu���]a�]O��T��Ϋ�gQ_�`�w�k�]�R�R=�Q�nCu�f��/ܴ����~��)Mوm���}�o9�i�Ș�_���T�i���� J�5�H�o[��K����;�`A������{2Xa��ZT�W�|B����[�i��EH �~
^���%�WX�JBs�2,qe����xp���<�;��p'�ӳȁ�$��aQ�ҝ>�$����.�f����/-nV+�_��!i�r��Y
��^(�y-�4����S9.�lu��`c���f�uḈ#��W�ơ���0�t�R��M��#���leOE��9ȳot�ی޺�ˣxk����dF�o�䀀K�8K��4/�u�ɟa��Ue����1o��mK��@�7�aƋ��f��2�_=��\L����F�����1��/��9��Gc.Y�va���yݵ=���~��e�]�h�D�M/0���s�¿�ȯ��ȭ���uaDu���@6������g�T����8s�CY1l��R�L�	N�/%z��-MwOC8�g�;O��& 5K#��n��ID0��]��G=�v���HK��y�ߘ�||�"z����a�$�ckġ����>�o���]�bR �(ga{&��|� #�z�G�N�8��bƤca�K���C����誕�eok3�hƮ���k��G�a'�,F��4_ �b�UX ��Z �Kp���0�R[����p+�WH2�&�mR[�>u�#�l�Zk4M��?+�Y���I�)T*X�;�-T���qu�U���VD�Ѵ��gL^���jN:����*-xz7�?7ʧ*�@��?A�QQ�ܑ0��L|X+�HH�Q�����k'o��?���7 A��-��{5o��8��z�}�8@I���f��,��ɕ�׼�=J����Z�_��C�B�^:��?���fL�$��@�7<��钒Y��T a�eZ�+D��R�&�yW��A�]��}貕cQ�	�xK{aq =�u
-�����a'�,�p):j7��}V�|��T��z�.�`k��G
2$Y?K�󱶯�F��7������oh4m��{YRN;��I�k����`�F$~�A����<zS���ޟ�a�k�`�w7V eb����*5�B��l�p� �N�,
�{�X���))w�Bvp�F[4n�8�N[af��k�+�qEEr���.D������,�_�t��Tx�ҩ�� ���+9b8T����F����d�M0��D���Zù΍�Y���q/�(�/�)?2\}6d
LӢ��6{���z2\�K�:���K���
��,r�A+�����G#�D1 Usܔ�'�®.rb�NVO�3�U���7.z������F.��`�mxWX��PQ�b�5.2.Z��빕�sA��&;��O�ꪳӯ��%1��/���.)@ٿ�M�F�ã�(��7� ��5o�zǃ5���J͆r�2�ݐI��^i%D�)�ǯ:�a�q��M(}��&�<���M�`d>�P7�Lp�	"���<��d�o�v�s���-?ͼ�ys�T��c��c��B��Y�W�"�?_�x�ޟ��D�ؚ%�9i�d\������ЏհHlw�W�P^c�kr��Y����-�n�8ØQ���?
�I�?�K�62�	�� _H�f ��c��D��<�jG4G�0�Y��E,�Ǚy�m�ԨK�f�P���?�ˊ+wK���6�)S��Kc�l��b"�����H�B��ǃd��T_}Yۃ��ؓO������
[D�O���k�[a�۩�aK$�����K���?$�}\���-I��ٞc
�ӄ
�pĩ1'=B҂a5�O��#E���w�h!�^A�=�*tW�U97�̔�"�|�Gi���j���zR�s#���B�����f�G�-�`�U8��N�d�3�i])�8����F hp���Wó'N�&�nk$���:��3f�ޡ����_�J�XA�a{#˴JJe^y�r�-�y9������(;<��;脶"̉q*b��J$ݤ�E��I�i�,2��	�y4�
�f(-���Q����ؖ:�������+X�׎a�e�$S��?�XL2�󦟞`�g���`;�7L`��L
�Ǫ�	s4Wl�������U6��Y�4���L|�	M�9v~q`�,�s7�`r� b��o}6���#)m�g�L�gW�0j�e��#����| ���X��@��:�s~����9C7��ʵ���&�<���!C,��@��T�$b�.�2�@��;�TΙ�O��F@��F��X~�)�vF�>r���]Wq";��-6#��]�GQwΫ���v�#i��c�(��ET,����#�Q�$Q1�U�0ˉ������B.>��U�����\�@���?�ގ���	���@8��	��+h(	H�FR��)sXMt=�l�-8B�Jďm�Y��?�X+�xE\&�����Xi����Q�� ��U��{�g&BE�$q��Z�B@��2��?�N�� �"l3�;��i�k�~,@�4����?�޲ ��4�ˣ8J#���e��t�J$���[�9Y��O�OY�El4(g��p�tSK��լQ�O�c��tH	Q�_򏿾���c�R�k��63'<m�t�p�I�ۦ�m
2)���@�P�6�퓩H��^$�H� ����|v�+ӑ�8c���	�H��?����u*��~{)j|z�0����F�8>'���P$Y�w��k��k<��1Uop3�9I�3���˨ы�]�rh+"��ڪ��$����-`�M��^IG0����wܧ�{��ģah�V֬sL��m4�J>#�mt/4�&����&BmO�%�H4\��'��Ν�5�ꙛG��p�;/�b�V0����/T�Q����L,�~XF�kB��i���;��W2����e%�t�ċy��Ĩ�B�ؕ ��.v�1 ������B?0���P	ͲM�$^��S)��n��͋�lx�)Ƞ��6���]�)X��2��B��,���ލ�B�ɝ_@$ihD��0&"������|�<��q�V3� S*�e�|��|�R�6^�g����-�������R;�������ߥ'yF�-ώ4I=��JH������5���G�.pܛ�*\�x0��z�-��K��1*HJ�BP�Ó�4�`΃c�5�;��J�B��UЊi�y��g�
��=������Í ���~�6�u��3�(4�c'