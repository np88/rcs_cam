XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����T}Hk[����֢��V��>̘2_<�;�&3�yY��q�M���c�����*,�u��5�H���*l����^�lSZ�CA��Mix6/��s9��PA�ت���[�L���՟�9�wz�u8�>qu͍A����K���]�6f�y�����h�ȿ�[?�ŅO�eXI�dD&��bqy81�]���٫�As�s��
��v�H��+�3��W_E�aݓ���N�A��5W�ku�,;��izpf�K݆����i�J둢�i�X��s4�d��)���'Ⱦ�B��G�(/+�צ	yc�O	�<!t=�`�Z�1Я��(��t��4^�zw���2я��#~���r�G���R��!�����KMԌ�W���ӑI��9�c�ggm���)4�e�F�L2i�fl�����_�Pja��On�A8��;��
tCr9��z_c�-U����L��:i��bOn��&�a4H^��y��Ac=9�_ZM]D�%�+����_�X�$�Oq�h��M�i_�%-��^�7r|��;�B&�Ѹ�5o_z�:s�+Xi�Hr�?g��X��8���$Cl�C1��N��1J���=͐�Uu[�������L�"`~�H�׸��bsac�ٚ��+��$L�:�6�a����sې�hjYx�c���aQc7_��6A�rK���@�~{�f͌����$7�����@��z�O�2&��չ�]�  b:����4�i~��T��8���&}�XlxVHYEB    fa00    2230
��Q��o�i֟���
|,�7�F:1 �aqV�0�a�Ze��[�]�ر��g��L�����%��>G��f�&�S#��!B�W
�i%�]�OS�߭cTV�������0{�C]^ �B�O4���OQG�;0ܸ�ugy���7�Z2����EZ��V5�αԈ�u`L���#�y�1�n�:�.�{�`Q����LD���G�')+��0w+H^�Mq%�c��!D1�(� y]Ӫ8�rd�^s���d��+���;�(���{"�겿9��6�@G	��>t�%p�Օ4����Mp���踱�"�]���f+f�h�ǖeH��¼��&�h�zE���S!q3.;H�S�����`A-�Wp���YbӕR�׽2{���i��(�)�u����>/;��u���fL�P�dXFkQ� g�E�w�5m8JL��t�_ar����ݏ9�u�PF�1=7���6���c:-k**����[)��.M�i=ҥ�g	WWb6�@��0yjtI��� �'[���!ԓ�_.Y'�]�ƍ�������� Ui�{�D'�U*�+6=I��h,c.���4a���R��ͯ[͏d��,�Utj��L��#���5Ę�b�;y�2��-���D �������FaS��ت46��tA��W�����t��<�UR-m��K�����i���oܪ��[��/�t����1���;��$n����s�J��C�J�]|�ݜ����[�����:eD����B(ks�)���X�2��@2�ۚ�|�^��-%у�ѯ���7fZE_�AEl^��A���AB���+%����cy��0��q]��Uxk��A�y�Iu*;��}���tl�˜�O8�mF�:�Z�ltѰqi�I�o�q$�E�4�#�ѓU�F��[�<�@���=�Y{wW��w��;����\�J��^	����UkI��k�ż�4��}�Ɍ�Ih]t��膋b韩}n
�ـ1�����^7p-�b����|�u����W����P�҆��}j�l��mY �"&�Q	�,${�>ie�een|�qSm�`�;��� �
��n��w�5$@���u����3`�R��F-d�yT͸�{Q��@#����xj�2�.;����P��.���kck�'/T��b�(��/�4b��n���P�}1r�,;��E�炋�ʯ�W��l�`aL4T��J�!�ɞ���n�|��rE����w(���X���In��Bs��ByV�:`"œU�Lښ�<R[�����YQ%a.�<?Vlt�bg������nQ�n!d�9�R��J�Ũ_����R���+yOA��Fj)gq|B��m��m�S�'0t`<-7�#/!	/�<��α=��	���枛;BJ6u�/F�&nC��G��H�1��ix&Af̅zsW �3����أ~r^� [g�AR�ޱ��Q}��~�G"܍
X��bL��Ґ���� ?��O6��+e'� L-��FS���~JZW�w�\��a䧚�ïc̃��0؝��(_�$w���R\S��{�"��1�%�0ӷ�`��L���+�Q�m�c_X�y<d�;���;j�1T���U��e��R��Ds,~Mp��b�pK
��wo�7�#R� ��VD���¿��A�WJsa9f�oz�&��M�ec��ڦ��2xU(�o��d~3��6Gq6 Zq��2��Z�U�>�����9��B�~5`H�:V[� �'��(�)��t������_�7w���S���T7Hӹ���M���6�H`tӥ>�hm��.�=�6��W�s����&�D_$�YFazѪi~��0^+(X�Ұ������5�S s.E��+\in�ƾ�;�@�����C�~ʓph&ƺ%i��:#h��!G�B���o��c�L�T���&��%��:�.j�]����.�m�|a���E|7�n5�M��ƌ����D˝��9r��,�e�~��9���})n�R�2�E���_!5��h��f��q��5�fF
CRH��e >:�#����1��vR:a��;�g��SVI*y���]�.[�]���A��䡰�C(T-￶C��aa$��ػyl���S��UT꿼�������Z�$h"��j��M��v��R4Z��_�Ɯ�N�T}=����LF6�״��s''{~�`�}�X���ҥ�e���	 d�N}���+?QwK�A/�/`K���3H���j5z�Rp2�3��M~q��۲n��_�ư�ɷ�oE�F�X�ԣl�J�I�'p��^���tԕ;�.\��ْ��'X��G5��: ز��A�-����1�7�i;��	+�����k
eT*�(��'
�*���k�L���=g�1���[�Q����{A��_P��XC�j���]^?d�K�pWb�ڍ��`d����-���E瘭pҼ�QpaK���5��orR��]�*����O��j-	>��9��/a�q������5OL�����琀���2���u�܉�n�,v�@���%D�s9�YJ�G�����s�~dm���E����FT ��D��G$x��R�ԋ#��N�+��>S����L��s���W՛멑Xs�zPjD��6�<�ߢv˖���������ߟU%4������8�|i�>�У<\_�rc�`�bV7�����V�����;�˦T7{���d�Y�/)��9tҥ#���+��q��P�W�/���-����7�g��R��w�W�f)Ӛ�mC����!�=���:�a�?�ݡ�룇�����W���N�I� ��i���| �?;�/Nc�8K;>^��ܣ�t�ԇ��=[�]�f��nPBh�P�w���+���h~��	�5�gx��E��w�q���څJ���O1؜�����������6h��+�U�-�a%9�p��h��M)��+�Rx�"z53{�X���t�'�V��K�f��6F?���HB����zK�9 ����^��hS=Y�V+@沖K�}e���a�>JY�9	����O8���L������|;�@�Rq����C#��Q��࿎N"� f��)|�1��f^��>�O0�E�''@�܎��|�S���i+�8z���MvFA�T���R�ጏ.�6t�CWQ�P�L(<ʌH@��=^	o��Ot���*��E�A\�Ձ����0�$1�q�\hr
�X͕/����R8%Cݘ��$��\֎&Ւٰ�S~�H��xP��û���I�A���̣��F�[��3fi(��FP!�4��6�w-���;扯����W��}�`)T%��4�:Y��_:�x�B; �|N�ڡo����m���q%�Ðr�W��Xb#���iBLQ�:��a�*b�ƣ�B���(wO�ޫ,�S
�Vݎ��u�ذ\�y��0��|���ߝL�TS_1�dk?�]�Y�Lеӡ�W�h:�0H)�i�\�C��Y�53!�!�a4>�>�����A�aB�#�i��t��kspS���e����iaս|r�ΐ���`�s��^⏈xn� >x�����A���tv�[��Tg��`�cpνPJ�M�/׈��%�#	���>�K���h/ix��U�ս|�h�6�Z#c$9录�O��MMIzT�A&$��A�
�YhM���C�ܞ�*�ot��e��	wH�́ ���&#v�T������X�`�&B��g��ܺ�0v�l�������ō��'k6M�o�BJL%�wc�f  �?S�$�!B��m�Qs�ym�xx��Q'˂�&�� ��%C��Z��!j��qiuАsBN�e�V�Uv����P�+�&�����hqP��ݳAE��z���Ρ���KjN7��Bȝ"���F�<�m�e3���h��-Lx<g]A{'��fۙ�W��F��y���ak�B+��^
<��QդqH37�>x���Z8|�-3`��:*I�,i<D�sB��K7�B��:��.��lA�+�p�� m*�4g�@~	����r��~�T���!\l���+�6��Y.��ݿ����"^�2��G��@߹w��,=�{o������a�T��_��g!�HW/W��+�lg[��i?q�H�����ƨ)�F�8���~������o����J1T<vp�J�b4,Q_!�����N}��>*���e��;u�h��e?�ġn�;��f�$�E�AK���n����uҰ���	�y���J=����$}} ��s_�F��5�����o���Qj����$�V��'��?��T=+S��!v2�3$ƨ�����5(�L�y��/�X�G?�2\C��Ц��<lTF�����_�$�{9
�n0�S����-� ��."��I�����J<mw�%���{t�0��%����?�G_!(AFb���X�@F�?���2[OW|�j,x��[=0!ۉ�̼������� �+x��Q,�E��|2��?�p��HBF�{�>��7��n5@����u�%�1�*JU,�O���.6��,d��R�������}-j��;5EUI�[JK���t�u�x�:�:O�va���W�	��g���9�q+ <�6+H�*��"0߫a0��)�(��Ԣ�īW�LFr0���D8�ʴp��LG��B���|���ί�`w�Z<�����e�;���TI@�A=��l���E[��ĉ�1N��7׹zb>~��J��5;�=�	��=R�@���>����h�04� ��aRh��26��C���&����miG�q:�ѯQ���	U����A�'�A2� ����aJd�����KT�D�t�r�:A�4�n�?�<���OT7B�ѷ 𕤃Ӭw������}��ٱ1�����/�������>} ����A"��T��
JȊ���U���(R@�3���w���1�3$?�!�*y�%f�p�s�}@{���'�ύ�G�>��� ]��Z�ѷ����L2Ԋ;yJ뷰�P=�έ���Nj<����zAG�w<@�@�h%�V�}*K�S�'z�S�kA��5|� M�Jp�"�]�B�����L��:�0�`?/�ԀFb��ʇI}I|�e��u/~��������ᣝ7��Q������t������f��:S��.�N���"��4XDI����`�����A�U�S�P1�G8v�*������H4*ww�]Rr��������� @ވ�����}�0k��ݚ]����7�2��w<F6�p)7 �@܁0:c�4���z����e!�C���;�P���s(���Oi��zb���V�kKY*��*�Y�c*g�i�~`SS��7~���D�q�5����'�z��� jp"�VR;���v���H�蓯0�xa?��4b�cz���0�������§ǃ'��GU�vE��VH����fקnQ��������Yo� �����u���w��~�E�@h~Ð!�@rV����JI��)�oF$�/��4��P�-l�|�l!d�3㤌RI�B����Y��T�9I��hC���߱���>�$d;.�x��#'i��qCs��*��#ʑ���b�^����wn\�m��Lc���!;ı{d�!�S�h��*�Y}�����
I��歅7����ߟWwc.���7�%q�+Z�����d��b"+����u.�ʲ��Y��^���b����8�%��}*�¹��@qi䑹4`R6O�"�%�"�,������� ���I8�D��
��q/<�4�A�>˩~[��[Bc�Mؚ�,l� q�\G�[���q��X�u���m��QPw_�����T5YnF�2�Il;��&�����[�}u���yy�G���U&V�>&4�z"%=[H���m��G~�])��%B��]�����Sb���BP5�in�	#>H>�|�&��g�D�@��0[p��)L�Z �42b&�C!�����[�"�ܬ��ݭ�Jaڠ6�qOlz�d$o��m�]�$�XHq�cB
��|����,�(�"c�B��W��T@���;z������G
/�uz���'��|��*�|h�s�|��|A�6&��xr�b>#�B��Ǧa��S��_�ww��Zcp�n[��E�him��-�9�aS`赌�R�z��Ee���ע?9�!�1B�#��b�A����xB��S���⺟��Ɵ��.Ҍ�bH���
�L��we���GO�ҿ�v���*#�o�:Q��q���痤J�$&��C�ƚ�(f����ت��
7�-^�-��p�U;���k��a����/��yi���k$g�t���K���g�}���H�v�x$�9�� ��#��*�)k��$E0;0��)X����a�j��|��!2�����
���ѐy<QS���]v/V�����H�S��	��hB&7dR��v�2?��VP�b����O��=��@y����b��1]�c�k
n����O���z[XL{%{�h-7�O� :�C���1�j �*���7?�7勺����?v���˕��o�$gz09W�)��@A�(�h{�0b����`0�$X��Oש��09������k�5�ަ��?nS��ɜ/T��	mm\���
�c������`��=TPm8A����-)��C;V/j��l
�h��_�ò�J�iʢ&8�Sg��v۾h��#V����-E�]�^��-�ϣoF�^�C.X�7�-jt5.زی%v(RrUԧ�w%�^�z�#><�ԓ�F�-h�ǘ��������Iw#�Iݖı�+�,��}�n����T4���o�|jjo[���*K��Jk�A��i��a������y/\�DXE������Ʉ��A��a����ֶ�(�I��G"sf�l��HP��S�����ֹ��Ē��z���ЛJ	�^�:7}�G�h&�4X����J����c�T�Ld2�O��8�k��� ��w'�R�(��●:���@�Y� �!x���i{�V�t�� @��#������?�9tVjIx�`2��ꯜ���6�h'Μ/򱞑��~���,&�عb�M&,�����[����"�)��YͨV>�[�ؗT����)�0��e�(i/=�.|n�Jk��Z��9�ٞ��؈�ü���q���U�����$J�=�y��k������FV˯gW`��,)�9~`;���2�^�U��}F�Խ�Ɲ)P�����({���H��'eF����^v��E8�"�7
�6 �-�=�.*���t���M]�I��N��P�F?�Х�yK5eMY<{��rB�8��g?2tec�� ���it���p�oocI��a��Е9��F��(.�V�,�z v�����D
�@A���8H����吵�^=.Py�"]DzV��j�č�wA`w*ZK�ئM���FB�߮�@v&�4�_��+�dL�mH|�-��P���j��#.a�ZZ�2��w��:�͈��tl��T�P�1H�M�#�����B����Л(��B{R�Y���!���ym��**��иŷ��Ls���U�j����&�m@SI�����<u�.뛠����k���1O�s�0_���]ᵔ��gD�*4n�֦�.��
�ЭAi%�e~��>m0/�oҢ���xZ5��N�7�����.����|��Q)���c�c�Х�'px�X����Q"�~;���zY��k$�S	g��>�Ν1��,R8x�H4�7y�6���O���O�zP���׶z�)����]ʭ�V]�39f�u�=&G�.���˟*�˯�< 6�4��&��?�tS	� ��=a�"��ڕ\h�y�=���Y�,ಓ�j�����ϐ���Z���V�
�,�[YV1�5>���]ɏ�Q��rS���~�H9�N�̮��P���2X��(�����w�A�Vj�p�a��{��k�Zx�('Q�c��]%q3��ݖ�	�˸�C9OtN�J�����L��Y����Բ�nZ�7�F�S�2u{�	�䦧��H 'Ȝ;�u�4�'P�/��b�3�Ǡ����"#������|ڢ���>[�%<��w��;p��X�q9r��~�K�lA���R�-9a"�,�3�ʊn8��~��&���e�?t��R}'?m䭩�G��ȇ?���tqA��^g[h�l ��tE���o*c0�.�u}�<Y���i���q� ���hg2ZA}�X�R��`DY9^�~>ܰDπ�6�i��-ER�\O�ӫ�7jB(
ii��g���:�M�~DJ������0Ц	�ƕ��z*}V)����C��d5�`I����zs�S�ƞ���~�m�&ث���i���#cr@R�ہ���I0*�q�G��vk/(55��7·���ɠ�ՐϪ)���<�?�rw�=��Q]��p�pS����.�d�ɐlE�K�:*�p�X�5��e�����U?��g ��0�D�~��4쀼
�,<�Z�t����M6YQ�;q�P�ePD�Ή��3z4�q��v�^��?b���<%�3���v�+�*͵�9����J|��>� �a5Ig��#v��l��Pq;�L3��IJv������C�u���Ă��C���T7'�S�*&��]C~d>tv��ZS�Z���<�o6�g����:x�~�FN���XlxVHYEB    6682     5d0�dxN�2۠���i�O��G��X>ri�#a�귟���.�&t�����/�LM0�^7�?��5���w���*�>�([�i}���&�ڲ��(�9�>���2^�2^.�{b��!`��j6���U�.���O;RT�ܔ�+� @�L��=�ڿA��.7�_ �?x�M�:�.%��	�6�Gv��g9.�S8=?oa�m�3v�ʽ�'�0�ZU;���>׮�1�ܾY��j����m�x�׬�
48h�%sS�ҭ���D�,%&��Oȑ���g"u���'d��%��>�nLf–`rT:ҧ�=Ĳ?��?Z�V([�x
q1 �g�>��b*52�4:Z�e�����jkNV^y��<c�C:-��7jhy���/kd���l���oI6�Ui�=]�5����¬�y����[�WK�7gG�+����v��D�/d��*�:���:!�3#��4ҚD������"�Yy�i��g�hL�$y���v�g��{�r	�M�w��]��u8Q������e�n��@Ju �E�W��"w��c���#�پ�<L��O�Ɯ��H�FWu��[j�WW%cbU�>V�8�y��
�q�#c�f7��֨�l�#��؏�HB�}��Mf+�7�dnt��[������>��`"~�JV  ]t;��q�Q�p�h��^��.�Ϡg�[ܮ�iO�6�@���)�f'�e�.�f�����Ԃx@���`q����3��X?=w~��>iD���fE<��vIN�%7���% d��x�ťye��w�sGa������r;����Y�r������D���e:�u����K�2X>fN/hl���3 L�4o�������������il�'�f�ԚX��h�<�<����F����T$Ю�r1~�9,fDka��f�T��`"��JuZ(�<��N@V'�d����#�W���s��� .�4�=��s�>gYށ�
�Ƒ%o!��'K���Ŋ� �{a�O�m�U�2M��KQ>'9�r鄂�� y}���Q���eg�����O��'H���4�5?�{ӛh:����S�U�DA��g�Z_���c�	wW2�oY��� �)}K�u��c����&
���U�����HB�e�����ovi��SG�q�0N�Җ�߆@�@���y�g��9KK���z/��v3Y�Fv��&��ېa3(���oS��4g�H���t�d�5��F��
����%�	������AD#,-[�M!��k%�J绖�(8Oɴ�t��Ґ��o}".�p���$����D ]���Q!H��N,��ƗU�ڴ+mo+�����d���ϝ)��w�F��K9
�7� Vi�
-��}�>�ϫ�O���[����x��Q���1�\�%�"b�� �A�Xw���oÒ_r��!d�Έ���B!G���A�;*,EfPc��}�%�B�