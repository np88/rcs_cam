XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����$����z�W�I(O8��T	��	��A�<̌L��U �3q�V��5D��us���/�|�P�pJ[�ܜZ��Ë��!D�ժ�_�$��R�T^D%U:1��}��f�Rt���1*.�ڱ���T�N��C�qS��.k�Q�Tೊ=�nױ�=�dC=3Ҭ�����-ccyy۳J"��&P����Z2B��(m�ƪ��| &�'�o��|�he]��N�ü�vm��X!��l��2z0l�+kj.�+��W�>�`F�1���9<��F�I�k��X�)��Gӫ�'��D[1�e\RN}!
_��L$ጙs�K�0�	���O�t���:����Ր���b�	���T�\%���{ż����^ f����g��P�`���n!�NcbU���14�iw��Pb���5�Il������ٚ
�� D��
��.E���U��Ժ�4`l�4��S��lsSt����B�-��c����zRJ2�⣡�N^�]vb��d�O2��s��ע��`�:�ơ�q��|�j��i�R��z7��*U1!A����?EJ���?�;�M=�ú����{ �� ӈԪlO�\�8#eb��?��;w�rs9�^�{��|��_��a����j_7�o������Bx����3_�y u6>�U`쨲Լg?��Ӊ�T�A�Ȟ����q���H0�=gn5\sO��}�D�;�2헓�	ou����x5� Z�|�_�*��|��8�0���t��P(p�>R�WysY��XlxVHYEB    6cf0    1960'zV.�!�������"=.O@��=�z����L���w��[~�[F,'������:b���'��@�QO,L7}��JR��� 5^� �@|�I��uhlel�
f�T�w�o7�V�-�2�L3Kޘǚ�]�/��պ�<N`������kuv(Ҋ�F��'V]��yK�^N�������F����M���bs����j��i���A�s�ݦ��K�Z��)��vx{���Vѓv�g<a!>���}�4}Ћp���$�t�E�{Г��.tU/����gX-+�w}�hk�~D����ٍ*8B��EÀ��~Ξ�
�
���Z �h��z1ݯ\�YW6��fuL������xb�t(�\9����Q��;�ԃ���)�ܣ�g��S�����E��U���ץK�o�%v*���e�Ɋ ��'M���d�G8Y��u/!�w������pi��
co<!5g���f㪝�����$RU��^[�nEZ6 �^�g�8	��4*@�*׳���8�������1�/�a�q"�k�6�QՁ��dS�^9�YL�d&��(3�V*��0�/RO#DA&�8�CW�\��٭M��嫊��H�S�_�t�졇��Xg����ΐ�]?�<Y��U^:Z�E�{�>��)Vc��/��W'�u?��R=�Y�Z�$��u��������YJk�q���u�� ���B�㔣����l�^����y��H�Y��x��Ⱥ	='/j� ]
D��u�N���Bo
i�So��c[s����}0�.g�BM(��P, ��:
A,4�BL�Rts�ng��@fts��~-��]�A/KB�)�Qm�|@� ]{��tWx,5��odQ�f���qٜA�x�����ʵT����	P����O��!v`�$����4��0sԵ��[�sZ�`a(YG�.���/��Hǫj0�X9�;/'�"��:+��*��"�6�j�Fr����x?���^:I�&iQg�2�V2�az6�<|�7B=cG��i�N�_�#io�Og��A�֗��M�����������-R$������i���C"Wu��a�=x��e^M��|Nؘ3zUQτ ���zQ�+�.n�
���9���"�sޏ2[��,�@�T�ͮB��/�[5������KpG�{���)�x���itz��^+�/�H֠��le����菳/�^��ge�:�j8 �T�j͕��D�So������lrRa�1B�ja7�x� rԆy�=z�z���K�!����(Ms7[B���i��O'�7�J�IoV��1�w��$^1��K�:٦@�r�3:��%/��9uE�&`xX�o쏫�зM����������A9�D%S_���l�͚����u�(�h�LxX�bmʕ9v'DK��5�5U�á�s&B���e�����ѵ��r"Gx�iֲה�ˡ�lSɉ�����`���H��9�w���ä��+���Xr���P=F�*��$[�]�]G\͟H�^#B�r�F8ݥȾX_>LC=�;6�N&ZB��yّR�\"�3V�*һ_�m[G�>ɫ������-�>_=x�ݮUx~ en��.���$���)!j�<�i�8d�~� �VK'O��y�ZҺc�m�49��GT�v����;�4d,�� ϔ�U���
���b���S��!�p:�Dұ���W�. ���0��K(���U��o�ܩ~�לTm-����+-Wj��6�P�vOt<KO�y؉�˹��;Sk���F -�et��y�ֿF�f�����"᫏i�B�.�ވ&//�Rd=���a���݃��6����JD��/�W�[��^
aY�J�W@�q��5�@Fni�s�݌0�!�X1l[�1�:Z���x�V63��Oe��p�iǣm�:˙��	k/���qR}͓,l���Z���-��}KA�GG!�<�1w����R�W�j}Ck�O"rqh£*h�@_�A�i�c��e�>��ঊM@[�n|���,��"Yc�|`އ�A����H������uR���lJT�j}�i/0:k�T5C�Fz��8h"�5����1�� @�?��=:.9���1�$#g&�y��TZ+o?r����[ /���Ğ]{� >�g��YjPGq�9�~k�Sv�Y��P���������<ݮ�u>�G���4���y�?��:���q��8^�Ŀ{��˩�������ԉ ��m���D.�OF4��XX'�3l�� ��oW (��}[��ăZj���x�����Rݳ,�#;�&
�<��d��ro��lmX���W�� �� �}3���/ �ɤ�*="U��C���@I~9�L�	�v��N��(W:�8<G�N,;��R���k����LsF���ހ�>��F�����/�+�l2���(�`����e5.����Hq�f�''(�|oA��;@���&.e�s��Y{���4��HA�p����I�S��0��G��Msb��q��f�6E]	
��["���7y���/�'E�pE��]}K�Ud6��� Ƃ�N�6k����g��
���"N����u1�k�Cl�`�d��<�b��z�T��gu�y��cӭ�Λ������xt,l�Me��a�g2�V�@�����wU�ZA������i.���;G���+�_���6p�j�B����Fn}�f�R�L�5��C3�T��Ð�=i4�_��(h����x$����x�9u��y85
F,��;A}�Ry��׫y���S��1̖�B�vf����p/D��)� ���X��%W7�[e�L ���l�Gq�,2�s�*y��nV<��;q�Q�)�(����j�LSi����a���Iſ��>�Qn{�"?�����|R�J�Ec1�\^ҟ)��b���Z'��\L�^���n���#���W��$�y� �5��"]��}'&z�^>�7^��;w�^��'ll��p�'�Í;�ؼȓ��Q���NF�;.�HM2n��?�O�'����݇�-�BapѶ8�>9�q����ǉm�s�塸p/�HW�w�5%�Y3��u��l[R5�ѿtZA�iO<�9H���F*���'9_Mn�Z��T�c�S��k�w@5I�Ne�f���� ޤd�sP�<x��GV7%q�Kt���<�]9�#��>��{B�b�O�^!��O0��84{��_��Je�zv�_��n�lM���k�m7p�I�Xs`���{
�}Z/�ڟ��-G��{L�M�6��Θ>�I��;�P���<�z�B���i�>�$F*��`��?�T��I�N��D�Į<qRl�'��i۪c�f+�JJLT�]�\�"�xd=5B��1&2��q�VV�8��N���_ N�x?_�h��{pmi���\��[��+��z%�w�GD�9�[�Q��tC�����;M��q�k�5I/'5�9����,wٹpg���Ca2%2�L;�>����R��j��F1hC6�H�\��r�6Ѧ���49h�k'��\���C��>)';�:�kY(;�po@9�%�g}�#H��z\�#���}�D�FF��8��4� ���[)U����J]L��a�~!�zߊ��iO��\ޯ���~[�)Y	�|����،�h�(|���D˂�3�^��s:�¤��2YH�ecw��_�Z�KӒ�s�_�ꈆMw�.��nvqW9-��ʠu�R<�Sw4�TNM6ܗ7&L�0�����ӳ���ewW�b�q��=�Im�Dٙ��|�=�*Y�`�� W���2�D��~a���ix�ĭ&5�$�� �Fa�^s��f�g��q�Z�cW,��
���o�uff�;�`�����[�.�I,���"��Ο^�5����|g�+�(Bf�~�|~��A�x?G��y��g5�޵��aF����u�(5��t^@�p m���BO���kɏ�Cޯ.ٍ϶
�A��;<Q�W�����?�ޟe�S`���k�{�j�� ����C����M��J��[���U�wQ�c#��N-���s�.۷�N����r��,��:uFHR\5̂O.:ߌ��@GI����R�Lr0E�	�K�������P �:=���#A��f�u�]n"�:B!�f�ذ�}A���p7���`�u���Ι'A����{�X��i�>#�`đ����a�Z�S�`��?�pFgq���HR��j�ON"��t�d�;rB�yu��Ds*�>M��D�w!���vk����c0�hxO+	����(�7����^lal���X)Y������3V��}Y8&���B��F#�5�tGꨝ�D��9�K#B0���;R�����0z�7_Q��c�Z���������Fj5��QD�?K�.�s*��iهh]"7$B�n\������Y�T����m�S��`ֻ��\Kh"3g	�����������z]��IΫft�W���J�B��{�8ek.�8>�"�NDz�B���=�SAB�O=n��01���=�B���נ=4�X�[��)��C��Pp���+�!J�������r�q�3�u��),[�1&�y-Fb0L�*��YȺd>W���+�*���q�i�ث�y./�h���[��'4���;Q�����ġ��͚尽L��3�@�^w跎�ʃNش�p�ܪw:
XW|K샐ß	��'��T�ҟ$�I�c�.��h�*<Ι���
j�I�U�?d�Ͷ�Q垭�5��x��y�ud�:S��%����:�uY6��=�.���]>�����M,����=sh04E�u��bBA�Ƕ��T3M�Q�$�ۋ�VzM��1�)�ˈ��U4����M5�����ѵ�cWM~�EӁ��:���C�	Rd��ڇ�w3�C�"tGэ����]_�g1���ά)�Jn�����Mn�� b?���"ɛ�)�ԫ]v�,��� x�PjI���?e_�ϣ��-�9���3�#�Q��W���*��l�]i�zn��L�~׆fS�L�������|���Z?��~t�� �6��<Ӥ�ӖY��Zi�����6͝x���t)�W�(�E3��¹8?պ~pť�(��B� 2��	��
��a&88>�{l/S
v�N���V+CiW�F%���x�9��#��tr$�h�k��r��Qn�s��N�����F�}�T��~�A�68V<�r��D����df/|�a���z��_�X����}�/Z�4�'�쓄!{�t�k�F���玃��&n_(��G�Ms�*�k���2��~�!~�Lvd�j���r�c�u�=������Pozm��>��5T"&@'/�fT݇ ��	&J~��GQ�`Җ�����G۽hL��$
�JȆv�f/�/�˾���s�?�檝_+���qGʌ}�=����h����Y����i�Js�<�E���Ǐ�Q��z֎%�qXϮz�"oBt��
3(�A�1�\C�'����[�h�WpoӞ����>�/��|<����g��xp���'Kȡ���1�r��нu�c�<��`�{�3��t�:7�0hѬX�c�����nx��A�PF0�E��{�t	��X�i�'=� �O�9�U>H�Z|��q_��B���;���B�ܺ*\f<���Ko ^|[������lv~8�d �A���jz�H�-�x����E���Y���cu�{�S-r���Af�"�;��Kl7Q�ш2�4�R�c�����r��s��4��ﺧ@l_=$n�%���F։�ovT5%����Y��XԳ`�?�l����,�t�IV�����ύ�ȱ�z��H�|7�E��e9S ���Λ�\�O�ߝN��.b��V؛$��2Jey��"���E؁"7D聏��X��iI�Ppj@2C���ي�2��
F�/������JB�w�=��4�EQ����m� Χ�h�HOY���
��
^Rz{�C~.�Ta�ag���sܡO��D��l�Qn�TU=��j�H������n�J��c5�1�&m5���JL����HW̲����R%��(	V���E��=c����S��Dٝ8S1+k�
�2�+T����h;����Ԍ5���
1lC���x.�O4<�U.�=��=�n�s�3`�3��G������t�kbY�����V���j�x�w�,uKzG��3�wk�ѿi�����
���(��dt~B�=U�z\���X״�krJe���������~�������Ϭ6T,wT�c'�n����`�?�����{#��kV���.]��2�-I����ȬAl��FG3�2��Ŗr�#���F�$�,�N�!���1.g�{P ���MT�U������
�t�?��#��+�y:@�fٜأC!k� �٨���N�P�DB���