XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Y�>��6~ú=:�z�^��M�2���5"��_�K�V�k��q��&
i!��k��&���a`>��Zcf��5��H!��?��m���TԬ)�J�]y*0��,f*�	q'��ƃ�������kX�/!�d�y���?��?�`Y/���4���a��Dw[�]���]��Tb��s �A0Y$^N��}ޥ�_Z��$ƀ�Ӣ�-��X���*8���W����;X�/���jq�[	bu�М[߬u��h�MR���Ih�2�(��KU�ܑ����<�O]�$�/X��F|��!�,�]scwWȊ��⚲��@��c�V�2�G���7�o���mꂦMH�̝,�67�ʱ���@�.߱�F��È�����c(F΀m�|Clu! �;��S
�|��~@7��YS�\��n'0\cq~�V��vt��[&��B�3z��  �~^�}��];:�6'{t��#4��F�@�������,�v��9��U�H�F���e�+^������4UR+����l��ۍV#�y���G:Հ�Ǎ����D���?���D~� j�6�i��vzV����0��3�3�Ya��!��N&�ظ�(��w%�3�<W�;q����g�WCQ�;����8�5�FV����$\琔*F�K�#<�����̻tr8~�Q���@�V9ʦ/��h8h:��P��𤸎� ����l[�~W��Od]����b?bO��%cgy�k���������kG'XlxVHYEB    1ffe     9b0���}�x#v�V�QΨE�ZR<ɻ�#a�8��� &^	�P� 뒷6ym�����^$�U�%[85��3{'�ͮ���N�α.���*�f��?a�i��=�s#�)YO��yƁ�qU{�X�E �Iҵi3���6,��ǬT�.�'�1Z�/5�(�A���i׳Sr骼�p�~Om#�$	�� *��~�/�F\�OoM��iє?���[Z�V�<�����>�v�7Y����u�nF�Y�g�k�)Cӻ'B%;�t.�=7�C��2_IO�t�<.�e���fܮxF���;���6ÝW�"�7#s�҅�ɾ��ͽ��%+KgD�^����AU�$���m��a��;D#J�T3�/�f�TNR���6Ƥ
�חZn@˶ ��^��AtIm �6�T� �$�@���h$is�T�$�4{n[��6���ad�c+�]�Ls�$@��h��r<D$�Hq+����g9� �Ą:pl�yN̶o�g��{����)�(I kS�`�i�FP����@;�P�>}�0dM���?:s/_��K7�f���Xq��_�t������ؕd�L�1��-���n��,eIU� �����N6�+�b���i7L�3�V�ę�m.L�`?�E�tg�U����f�O�]rb��%S�Q?��u�<iO�Z�Vj���^�3��]6f�p��^��TT�����q:��8(��-y�Z%L=&�܂��e8h�O���W��j�?=�=$�Wh��D�=	/>ڸgixS5��Ug���3��GW��	����s.��m:�`u}C{nX?�\՟��@a`�=]ֻp�]��C`�f�	%W>�N��S�e�K(�Jo �G�g�c;�e�M����MM\�T��4��5��I�r��Y�v���'�Ġ��ɧ/A���S�����$ĖŴ�C?�c5��C�䨺��pj��ze]�T"���2C!�cg"\YI�w�\��%���5�t`UO�m�(��A}J�
=�#p��K�ygV�D���z>	��$�
0B���%��8q�ZT�~��XHp��W�1%���D^r����������HW�7<�)Qc��ߧ��Μ��(�׈])��+iI��Hiܒ��T�����϶>�g/�����}��jd?�����浈��TY7��??�&H[5�v��h:r2�	Ѹ��t�� P�?t������ƹO�}?Ow`FK�O�H|��-[W�����s�,�Muz>��:2"��/����¸��e���H��3�Y�;���,��ڛ pl$a�3��|�E��/�%��G��M������=���S�7;�/nx�+PgA&цܣ��D*m~��9?�n|�#b�t 5s���/k�Pf�4\��9�Vr}��i	@Z��0����F��2x�V��3��� <[Q�9,�߉:��A_O�l�`�G�E�u���T�E6?f�����4�Sd>S�g(�gF��L���P�Wr	¹���l?e�(��`�f�
�T�!#K�*yą�!op@�"pH�[={-���ȼ��w8gF`V�����D��Ma&�K|��7�ς�R��`���U��� H�T�QE����g,��swxU`�����$X�r�������<�>�v��nh�����qK��	��|�Ђ��	޶�ib8~�:q�v������7�	@��7��g�͡�__�<��T�F�ք�^�B�P;�4��åy+�3Nആz=(�k�qi�KKP����4a��҃���Y�����*�i��8���W��ݭ���J�nCGM�x�����_[&߇h}R�܏��\�0k�������a|ǈLG�E�֨���F��`r�C��̺���g��I��X+Jf�K�<�Ӛ}ŸC���+V[���۱�t.�2�^�u��H:33m��/���񧉊:�s�<Y��H��B���=��v�k�c�@��F
����m�.��$��^�t����'�w
;��'�S#X*�t�6ͪy��2/2m��F&'���Y����O�L5�J��J�&ai���F� Z���x�-<�(pmɠ$�KX.�О�ܨ�b_
o5�U~��z�ДP9Ŭ�
���.�]%�MVPb�
�/�Q/�u.�=�P�l'����D����^�^xg�uӱ����$�$ic�����6�# +a1 d��I0q�N���5K�.=%�G�<S��q���E���Y��g$](�����;������"�K*뱞��	�<Cii+�7t;�/�ܜlQp�L�QtĿ���zT�d觺���.�EXeK���.6�(D�_�D�P-��εQ��6���\�N~ϸ�&
#�8���-L��fｷ*FJw�q�`g^Ql�-5C�[�f�J��� ~�DL1'�$�ex��U��ڢ3L6������Fo4 ?px���T؈�y���kW6q�N�W��6�_G�8�@��G�ˮQ��m��W��F&/�����}��