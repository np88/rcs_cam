XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��������-f��ѣ���f �6?�;6l���n\���9�����q�c���Stk*���C5Sf��8������{�6��S��^�Q�g��C^��ǆQ��v_�3�AW���I�F�q������)W�2��^��BP~�x���0��P��`������ivx��Y(�z\,9�"O�}aL$Eg�,g���#4 p�y���.:�d!����0OB��s�C0�� ʘJ�Z�g�}o��lN�UA��8'�?�����	��JBd9�|��q,2��>wG���"[���o�@��.;WPG���y�(��F��:�w�<��(�VC�ūK�i���%sg��N�?����"Q`�2yc4m젊B�P�aa�At��W\�R�Jk�d�a��B��\��ҟ��J��W69���oh�ܸ�	�=�.�I�������&�p Al>7���f�bM�|��=N�t�J�ؿ���j�[Ҫ��6��:��(²��:�#?�0.&yϠY��[ɳ=A�a��>�wʢ��]a3�a��ۧ¡�u��Dt�q{[� X�X����\�Ki��v�؋�̑Y�Έ���xN������㧏��z�/+��V=����6�W�B󽒍�` S�?m�t��܊�\à3V���<D�cbF��%�B�A?y�*uQ24���u:�%aڔ�v�D���Z�9t<���A�u�e�e�&945L'qe~  �.�J>�7�f�{�Ԕ�ϻ;�O��B��B ���Vt]K��O�c��*���D�XlxVHYEB    4cfe     dc0{�w?�1E<��h2v
Y�J����k;��G'/�,�gqI��� ~�Wk�����z���Z������E4	G/��vkF�H!d��H}B�u����"��ML%�A�vd>&��>1��q�p�q���~5^	`�5�[K��'[����$�+�ͨ�A��Z-�u�� �����-�vt��:@e�y��7 pf�.����$3O_m����q��\��ʴHu��r����c��o2��*�@\s���2�ě�!S8"�
6D�ɰ:�Lu��m�]f��,��Y��F�Q�V7���5�ՊiT��~F�'ՏM�LߘkD�W;,@�K��p?6ߜ^[�;X�6��/���Lڟ5��P�S���y3{0��j(��h��C���*�����������}&�1Z�%�� ������@D+I�g OH�I�b�Rs�`F�������Xw3כ�s#+� P��kl��Cx�hښ]TǮ�G �FX�g�{
�\�pwM�2�j�7���9�q�q"��������˓�D��>�]Qg�+I�j�.�Ky��Zf+4c23L�X�C��û�۞!�q��(���#Q���Z�T���g�r�isy���D��^��L:W�3l�����a���[���V� _�>��U�a8�k�%�D���8�&8F�14�ӧp��K_�ϡN8��n�g� fC�6���L{ixR.b|��}%�q/H�_�8�{�Ul���"dW�����3�{�V��
s�ޗ�e��ҋ>{ *`�#$����k���3�. ;�����Zn�v&\��z=%eKǮ�|ئ��n>FF� ^Dqr"=�e���ِE�����l�(إ��R7_aS��kR4���#���1�gZ${/i�di$��O�8p��<BJv�)��p%��V!���ש���D�1JfҚ���.�8���p3��^y����!�ynsr��̨鍼[�	J@�&�԰?}P��x����I����g�C;5�yd���ɣq%�3��М���X.?}�qӡ�FQ�G��C+ʛ���3]@�ʪ�Ę�y������~I�B���M�\-��-M�qL�o�R�4�������w�f�Pd��
N2l*����v�L�<ĝ��
�K���d������>D�c�lp�����:W�z�\�Z�y���HZ�XP��X�\"g�H�:C�{��~1�*`@��ek�P"'�����W��)��n{�?����|n�[	�dAa]X���7�����!]�]��ʂ���d jF>-�X�B[$�O����C�7,�>�Q��(����"chr���#=���ڞވ_L���!���F��A���rI�`rP��������;�DRHOBS���8��!G��b_�R6��T`V����/�����##�bp�>�R��ǻ3��vί1	A����1%Ŋ��N~�raܿ�v�ࢷ?iX�e�=���2�{￤m����Μ�kG��ʪj�T�6�Nkc��r ����S\�~畽e|��~w�$�4��ܵvch� ��NaJR���]��vkL��:ІeV�n>�-(VZ���Ȑ$�C�ED��1�~0l'w�e�e�ƿ�N�&��p5�L���gf��UY��2���n-�D�z3�՟�1��7'�xz0���\}|�^�P'�-a�B�=�V��J2����!Y�[����拔�����"Oc�U �K���)ӊS��YU$��N׏��Σe��
W���w����c;z��;�F��+�����o��N�A�(ְ�}�t�E�@��l�>����j����+��<W�c���&��4g���y��_�eYP���J��`.�b���'+�O<g��T���J}Nf��b	 fQ�I`{N��jҼ'=�[���q�Qm����0���$h�d�]�����^�L>�5bq�4�,�[�CV�ş�'��k�wZ�bD���ݲ��<�D.^j���Qa-�k�uU�U���C��`
��֖��!y<�9YWZ�*�[) ���50��[dg;V\0G�n���zu�����%�?=��^~^��+�**z)N��Zx���b}_��Z/>�^g�����B�:�f��nE�~���r�-��\�e�a��<�B��W��6�H�� �ӏZY����UU�J��,�X���]_'A!nt}Q ��vҼ�e��F������J%n ���תU�$��x�fv���a*�I?�)�by��.E�c+�(��Ⱥ;�2\^��X���ٛe��	��&�_��|��У���1c<R�9���n����t���/*v�dL����d�j�v(���D�c�$�a�V��28*X�=9F<� �-��ߛ&�0ճn��e�8	��"��j��q6��sU����� �%)�3~������܁E��g��:F�5�<�b��,�F�ÔO��T�h����že�
��CՖ��Bz,n,j�&0�7;����YL^Jd�B΄�R�4�'(HM!D�����_��QXyC�<+����//�I���GU��AI� m�M�
���s&n�Zg>�P>�ITn��Lc�p$2����������6�]�^�Ie�/�ɮ���l6�B9��lϚ.��9�z4���J��Z�Eo<�e{�E�Eu�4�N
�ܷ�F	Z�g[�b�����>�~����?[�6�1�Gkm��B-���܋�q+�Ll�nB�,�vW�ѱ7²=�\41 <�����(B���DY����͕��T��������z}���	���M֥H8�;�|�{B	ѧl�RMx>$���_�t]���>I���Ǉ���H���)t'|�T2Bj'�D�h����/�����2��X�'�CS��tOF+�k׿�n���ȷ��B���o�G?sY#�f��%Ԉm�c3d�����IN�)��M6�iB	M8E��,�2BPIGV��j��RE5�9~�/��3����ˎ��D���z��SV��� Kxu,�դ;��k�4bڋK�ƍ�|X���]����`���8u�lZ�l�A5�j�Ù�
��D�������q;�<��WTtTRg���R���ܦ���������š}��HTs������[Ś%|��Aϯ/��q��+1�v'�2�<��ߠJ�!=)�Z#���|�{�@Y�k���y�gR���0�d0�}lf��7�i�d`B�/��l{iu;��(^�XzM�~�Cm�5y�	ԭllϤ��1*~'�M�g �=jk����b+�kDn�lN�~V\�k���7����(��=dY#P�q`��S0�i��IL�� �~|9��MM��#��2�B�4&L�l���x/ܦ�2Gq2��y�������}ɢ1��!���>0u��}�����S�S�W�0��������ھ�<�)�O�9)���S		]W�z��!ews'��cvέA�ܜ���A������ �i�p�X�]ӔW��*�^���$�˱�F��IЄ̦�