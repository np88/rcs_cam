XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��/�M�1:䋘�"K#ihZ�	�)��w~?�t;��/���	�Ҭ��
���^� �=8B$�iBg�</,�z�L��{�M	gJv�F0q�����E��_[�fwz�"�a�-�O��x�(�-�&����K�1'?z�R�hH�.Z�����6��j�!1���m]���H|�FO[�����4S	@�oUi����F��Koɏl�炮�Ɂ��X�lS9b
Z��#�E���a�B	���YDI��5ƦH�!�Q��]�а��z��W;�B��Ͷ�^m����и��r�r��>�э�5�o�������v�lQ���i�d�o��7�':��'sOJ!�jA��*8/��)��_p�W�����l���_8l�Ȁ�j%[ɕM���@]٫��vQ�v��BT�m�H�Ҧ"S�o���������N�dś���G(������VM�)ې�oU84�5BT�M��LU'��x���`b&C�W6;v���Ҙ�׏9U���w3��������K"J�?b��1r.
l�5�n��`T�!n�4!A�$�hj�?\�t��=�*�62��;��������֟�B��d%ͤ���0~ �O��0g_����pރ�i���ú�L��]���#6�3͞�W[��3W������r���J���%��K\{�����'��4(�b!�n�\���Θ�bC�_?��d�g��.�(�[T&�[�x�����z�&(l	X����>��45q�XlxVHYEB    8990    1bc0B�lH���A�$��9ZI��џ�K�^�;�Q9˷��;�ݵ[�M[�KE��S���`_igP�-�@��0��-������I�^u����MZ��9",.��H�p���?W�	�^��
�=���]N-S8�c=-۔
���.1,d���[-��ض|Y=A&_��/a�Y7sY
�Ҩ����w�"�s~�ݢP�~$�z�BvC��̦o$ �����ϲ^t~�(�g�}��\X�}hWd���<Y���H�P�;R�t� �v(�K�K�}%c�_�Uy����m��iiU��)�jV���P�-@<D��kSw7�^Eg:R�r��	h21"IIw�yc?̠|3!�H������%F����6�K���A�]zI��,�� i%^�&��m�(o����醿~2)�Jz-���~C2P�u�hn蠘@��Q�Q ���f�����<� y� ���w�Rx� 0��/A����2�L���}W���T하rã�m��t�r����t}�?��E!$/��AO)����ی���Pn�#�+���ɰ��^�}��*B��	�Bz���ltt$�:˴��wC�ĳ^����6��
�Ֆ�Uu�?w���#Z���O:�Rf���^��z��7�g�"K5R(�[	8~��J��%��nyK����iӡI��x�%꽣�-�;?K� ��e����3d�&(x��I<[���0�&���������=��mbKx��*�Q���i ?��!;�H9~��zV ,�?���9���N��apǿD#W��~�x���%][$�����S1��V8�
��8�����r��CU�n��j��Pm|��X �����|����f��K$%S���r�r�G�W���h�� ��6�����v��^�k�lg���>��%<yug�ocё`�`�g����E�e�����mRi������@�
~#>�/;cI ����b��.�����T��?�� ��졜�CM��F��<a
?,n�������P9i7�ʵ&u��ؚ�ߧ��?��֖�ф��{Ψ[Q]:��s�k���S]�)�n��T�*(Y��"Z���]�/��EjY�,�����@��đ��I;��!�#4�lG�0������Z�iY����du4���q>R'.�V�i\8��=�Χ���&�<&��Oy%n]YeM�D�	��QSo���Vhg��79]#��c��Qc�0(~-C 29{3�-��J�eU�aC�����PG'H��#�����ǌ�Ϥ�Y��ĉ���w攬f?~�� ��4O�~�~�frZ:�F�e�x�Y�2�=$YHE\n����r��ex�Wb#�9+��D,6�!R��=p���kfU
���W�n���k�)z��#�h�ߝ�!�5u���j=܃3��'��p-�f��Tv�M&h��[�f��ױ ���	��j��.��I��u���g`��z�ĖH썁nO���:�K�А��0�'�ʵgN���biyFs��v' ���<����Mo��Q͏��c1X�s�_j&ȓKAC�S�$�FB��$� ��������@��~�n/��o0y�)̾��1Qv���i����*��^H��%-ɲ&��?�b���Z�j�O��,�Md$j�u��]�3Aح=-�'^�T��n)�.���1-τr8�\�Xa�1ex	���?:�i�JD���h��N�F:�*��ꅟA/�4U���i�M#kW�\T७�+!�V-��l=5��		Y�Պ/�Y`T%T=���m�U�s'�8*�	̧q?!�$I�}�`BҰ!���Mr4��ī�y0�q��*�`p�i`�U��)�g�y���^*��Ӫ�=2|Zd�9� i� >z1�3|h�Ade��FD�@���vH7��TXt�"jk�c��j��s(ǚ�^�R(dj��J	�8�_^5��5⿞�D�_�A�K6�b�;[�]w_9�3�l��Tq��T��"�&4+:$�'�6�tYA'[�B�9�5z�x��7o���g����}s��ˊ0o 90}yOCi:�H���M_��(��(b��5��3�,�,/@]���V�}ڌ;VY�� ]�dw8ݒz�P7Mޏ� �0-� 9�w��T �~@B�>o;�P�՝z��~L��CYH{��x�U�=B̥9����-e�򡻖��S�SL��<����+�V�J�:����#�7������Ј�ܓQ`�dKg��b�����O��xc���3��!s4�gba��:�j�e��Vy{-K�-�G-�=���l���0y����mLZ�@P��r�7�s6�b�p*�-����Jf\G�i9u��@�W����Gׁ��ء�W�I�y�UaWa�R��7�d	"� |�	vap�p���O�z7�mz�섐�Ca��ed��L%�3�)A;���r3:Y�T��GS,��H�YWw��I��=N`�^'�T���h`D����䄂�@#Q �S%�2D/����H�/��]@.@�)�n�{{��)�>1`w��GCd#L�����>Zv��2��Wi�����{�^�'��@��Hx�;i:�A��)�&���{�MqZ��$#@�|h!"T�ͼ_�
��ǌ>ޘȯ��R񲛤lop�Ͽn��"��M�~{\�YFho9��PR��+�D�F��.���+����W}%���Ub�ٶ6I�ڥcVL"���&����e�d���k@��>aψ������W5t"����:uU��H��lL��������],�����$��r��S�sf?(���x�����Qxo�a�3��2���<t�R���O�ih�9��O� )S����8�REc&S�� KIR��iT.��ia�$řs�?�ޚ�)n�ܳ��3���em��,]�)\7خB�u�:g�̆[v]��.�Y&W�f(��3�AR@�~���jr�_aۜe�T�=Cp]��Z�hΒHj�u���Ʀ�z��씯�<�ޜdYJ
����P��I��!�M�naB]~�Ji�N(v��;���&�Nr�4Aa,�]��TWɀ�@�:]��)!��a5�63J0[�
�~6��1V���K��(�A�K8N��,&�x� J\C��nFt������;���s�G��?Y����D�@�O+�t)�b#��M#�0���w�V�gi��	u}��qO,���-c��맻+��1[棠������J,�r�T�w�_�IGYi=xA�l����HC�
�BQ|�����w�*��Z��}p��6e� ��ȠYc��,�TC#�G����[W�ϴfB<sj��*�9���8����nB���ˡ]:?ݽL���w���kb|POX��uT<����Z��(2�5�]��NtV\/=e��x�=�䗌�xr��	b(��q�Jc����^d���ui�_4�6��c2�`[��x���-���GM2h����^RD0k�hT�f���&�Eӯ����I��T[!�����L���J%PɄ��/m-{Ґ��T��V�	i�P���8��,�3p��*G=���d˓<-�"ItK�8�g�x���s�e$#~�ǮmΙ��,5�	۰2���;��"�ŨμӜ�Yc�H)!��P�a���-G�0��Ƴ�=̡%������ˤmg����zP1���Α�v�II�{�
�1���L=_̮�"�ךA��A�}go�����}@V`�|�y�{��vy�:��ŞNܐ�t1ewċ�LKZ�+*���Z���S&��2;�9��;p��Q�j?|��ⓞ� 	`�������'�k�N�M����߇�y�a8�$s. ؗ�i��K��f.��f�W�[�x�o��ű��������b�m�&3F6:�0}�C�$v�Ex�k������rȉ��A���D��Ѡח��Y�;�DI�����O�p�f��(�e��5������;|�S���q����ţ�Ey��>�}��Agt�O��g7<[�+���z�����^�f�l��B���R���ޥ@٭!� TW���-����Ȼ[񇆑�y r��Xk�sD�2C�*�a���E��8�(i@@� 2�h�������R��X���{�O���`�D�H,��1�3����r��Z] K�\�0{#RDG�
S���Y+&���HI�X����tі� H�k��}�������~����J�#�"��������7�F<ZMd�{"�]0�=�_*%{`�����а�g_؏�C��4�쿇�%^(狇К[=(4݉���M�;�;ǃ�{��|?|��f]
�iV��۰j"W
k�k��1�XVp)��ٯ=g�1'ĵ����\i�e����%d�۷iN*�����ǅXm+l��'���׸0�d)?j/����ȗNK>�P��L�c�+E/�Δ�MźJ�|&\���7���{Qi\G�*/��qq���k�4�P9Ә$��3�y^�#�#�Ծ�9]��<�f9���@�/
9�Rg�<@*G��3oy�{������Y��%J��(��Y)�JT� ��N�W�*4M��,5�p��Q!��p욗U(,�a���h�N��ÜAN$N������fj��τ�.Ʈ~5.�ߨ|f��F*����Uj3?G��6�7����x�Y���wq{*�,5(�;$d��AInΚ��b�fi%���=ǃu=�d90N ��!��G,xLl>���#J>��^އ�(��>|��`���2�p�Tg��_�Zg��u�$P����Gb�P�ٺ4w��)ym4Ml*���*mu�9�J��A�[������ńB��.u�4�T�|�+(���N�OE̖�D�~*<p�ðL�D��rpk�,�1����� pl��ys�M�a�Z�h��������Ik��"� ��+�^�r(��&�?��R�C��m�7�Y��h�6�9@�IS)����k�Ԗ��Έ5,�ب۳�KD�s�)�pcF/2?4���U���`i�;�,�.��t�	րav�NF���pk��8[��.�?�аˡ�E�Q�ρ�2�Z�-�Krۜ^�/�k�-��k6{Ҍ�M��Y{�0*�����X��}���I��� �uo�Գ�]�>ƽy9�����p*9:x�?���SB�b���\�O�����-='K��9�)&�Bm��K^�hK?e�;A�L���xP73���g:�{�lkF��~9�¤��oG��7����ێ����9���r�ef�oi����՜1x�d߄n30�k�vs]�>8��?9�պ�O�x�y��8��"����!�vUQ9 tLI��"�&1��w��Yɡr�K���*x�x��u������%̊7�_�n���Q�Ȭ*�_�PC7����+�m�Y�D���҂Ɛд��dC���O洋x$���Q�W"��l�S�w�}X}yW�4�$��o�3��$�N pێ%��&u@�w������"�a~�`L~�x�zi��t�?K�[W���y#�M�73��񌯎�s5��Y&��Nc}57�� ��[��}QR�m�>p�2j�2��P{ٲ쾟��k+��XQ�[��=D%����)z�OP_����,�q��:lb����p5kOnM��� ��$ŝ#�?@����4�n��p�ʧ���J�e"�9]s�٭Q��7�T�0|�!�|���b���O7�����JA�%D�)W�\`�S�HX������s-4�/�kc�<.� �Yߊ��u	�8(����%o��C�� SPu�#�'�� +3�Y��@���]�B�M�d���K1n�6G�K5 ?DrN���Z2�е�^����=�$�j�}V�:�b�(f���q�+c���])}�qhb�4�����DB��]`%܉��5��8�d�y�m��Va��Ṙ_�q��\�-�߉�Z/w��Bj!m��)�c�3l��`��h���xY�ד�����u9n=c�o��5H��I�96ĩ�����Yf��~\{��q\/�䋜����vw�xw��m˓�J�Lh.�����x#������e�W��KU��t11��Jy��%�_jP"hS�B�DV*���p���ȁ����3�j� fM*�34�y�(���j��`z;b�Vn�T�@ݒ1�����=6_��ܿS 7y�I7ыO�@+�ks�Z
c��'9j,/+�"K�_L���w��#t�R��)�p����(�b��._m�}�?��7,���fT����z}���9�0���&q����d\;_P�&��"�겆ux��oW
6_�6�i��/�"lW���-)BX�.��lP[k��}�_BQ����LŅ,��ʔ�"bQgG V|� d��e{�}7�S��s��;�pG��@�lݬ 1"�Vf�e�pH)9lK�	afx�}�������� 7���3�B�����V�rt;%���R���>���zh�^��� I�G����@EGBW�.���W0�&o��h�a�����$�iQ�A&��F��+��[;G�1�٢Ĉ	B�N�Z�D��b�B�Ym�ܜ��e����׼�X��9/���Ϟ��ޫ <q�����*}j+�8<����9_퐕�={S���豗x����N>m�/�^~����}����ܦ���v������է~�j6����B�Bu1�1�~f�1$?�!�=�F�F*����f����#$F��^�)�}�Ф��<�Z�!�5iJ����씫���)ƹ/$CC��k�#�H�zIz�X��LԎtc�.��=�!W�����^��������"< ��!.��nY��˥��9[�c�b�j���81�gc7�&=�jZ8�Q�fz�Э��g�ص�<�!�%�$�W��?L�s�8�t:l�]%$Eegw2K�<o�}'��_?�5#��y\N�r�L���b�õ~5K�97آl��"�25@�*��
��|U�Z��5�q�Bj��16�ˋ�?7�&دI�d<���Nn@خ�;8�$I�W��GEP;