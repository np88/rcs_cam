XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��F,f\ �io��@����~��������d��du�����p��b�Mɇ��O$
N_+'G�)VDEM{\#8F�$5��Rq�Q�ᡰ+׭e�h|>�Ww8Bx����$�M�J7]Ő�E���`��m�Y*���Ɏ�R*��8����l1� �e�ؠ'6������7M�z��BtI���Q�1��������(^Y ¹s5�����ŽEE˃��: ���\C
(ʸJ��T��,5���A��P�u��*fH��X�ģ�0�/����z%�*`EG�A�6O7^8�rf1e�pf����e�ʽe���Hބ�p��zs�$	��|�r_����{S�9D\,��*@�N)�aL�T8���(��6�:��W?f�r��8�,Q��!w��\��=HV@�t��2��e�����{)@;ƅ��	Р�ҡ�z�T��]K�/S���O3��z�� ��Ɗh �)}p_�6R`���*\����B����Z�ܢ�vD��')%[�5����~	��,�����,�H�A�����}׭G�M��aFCUgBM�r��!x�� ��`����`=ki�)t������s��V�o�������W�]N�B�{`��̀!��v�*��p����.�*1��q���Nׇ��zc9O�`��#��L�m%���݇�*.+����Ks(Q��bYD�!�|Z �$
�;��U�Z@���%A���*F�31��,R�K<������D.|A�/���"��a�s�XlxVHYEB    6534    1400g3�%{��T�h_��&3�Y(��j,:S�c�Y悝��q�w����������T���H�� �f�(� ��6ᚧ�uQ�/3?�̟�z�H�^�����F�T	�:���&P��
���1���X��q��İ���a'�U�-���J��T�kƫ�]])�{.N�)fs���fJYπ'�S����a|2 ���XH���tÏSr�z#�("R���������0����yJ�<�U�e�}F�S-��HGoOD�����IB%A�Ěш�K�o
%�C,2!��$�5r�{~�p5��v-�J y�}6q8���Y�����s�u U�r}��Oy�S	���4a�RZ����?��.Oy*zv��WJ`����&y�B�:��0��k�?!?E���v�D����(��Q<*�S�*s�-H���O�5-?�3�>�F�9q�IŊ�s�b?�R�C���PP��;ѡzd�
�pc��3��d��E1���R���[U�S�O�j
�}a:,=�:�H�t�G�m�yߍ�j0�++�}�\@܆���{�A�e@�Q�.�T�]Gc���m���}�����A�
R4��+{�<�ӣ=���Kĺ��@`�3��U�Z�ۊ[P�N;�V����'=!��)b���e��u);�re�r�]�
��l�?G�!���Wm����,2Ok������z����_�5�_�q>��vy�s���dY�-e���K��"#) T�sZ���˼. �����_���u�,io#׫�V�Iހ�)Ҧ[8h�#�6۴p�1|�L����%�\a�*�!�8�#7Dr��44��U�
� ֮طڂ�t@P ΥIѱ�K
�_%��/n�+:]j�[W"��m�ۗ]'�B�u:ĸ��xLo��jY��$�G\%���eSP���c����,r�=
]�s��ǤA���[�$Y��?�ws�m����{X�P�L�-���+�D���V�#>f�4R�^�%D����Fa����Z���(�5X)Cb��I�B������0|�}�W��Z�W�9���܊~�߇��A�v)9@Ż�3���_������-n�	�s_c��w�"��;�<� �Ɵ�.����՞bl��a>,}1��D$����c�E�)�#!�&��"�;��Gk	�����4�;y��t�ȩiWR$/`�oX�{����]���[��h΄�0)=`�����W���X^8q+P�Y�.Y�e �{kcUa�tV�H��65��9�zH��0'~y딘��򔖕���{���G����:ޓ�izE���;��_?奤I�d0<�@ �^g��o7�X��\�]��U/;���������6�!�a�||Z\hG��lM�V%nTپ�ٷ�ɢ�)gw�zb�݁�sA���f�:�e��@vY���ZqUn�M,1aྑ�rɟ1�A���1е�m���,,��È�ר�eA�F�o+�t�����*-�l~��)r�����m7i㏘k��pe�)�R��Ê��s��i5���]	��Z��5���1���s�]�xD(/g�k���+�g1��X���i��	����<�z����D�F�4��X�ɽ՜N6����Mg`�u��+,�_�<>���o�le��ʠe�!����}\��s�����v�Z�:�	�5�àNW��c�W�l�iG�Eg�d�!�'�ҧԡ�Y�"!�ݦM4*!�����v[ }��!	q���z�xZs�X��Bs�N�(�"%�!ܥJQ�Rx�@gRX�$6���Kۄ����޼�'ӵǤ/ę�Ԕ�}9�`n��8���<&T��"�*c����;�y΋���h�3�\��O!O�N	����?K�ŢI�J��*��0`���pt�O\p��W,�}5F��ݫ��e��n��f�BtdP�昸 ���Pҏ2�@�&����ղ�a�g��Ew~���)���R��l
v'L��^�C⫭Z\��	t�Ыb�^����[��Y�`�ld��g��z�+>��n��頰�i%hn⮧��������Ҽ�����P��%�`d�c���8�ϧ�#B��^/����8Y=G������@�f�	0Mo�^h��q��|V���H j$��W7��u��`q	���RZ̙.�$|ʢ	�!|�!�iT��.̾H �h��%���,]q]��+	�@L�Z��n[��R�F����Y`���0�P@ �:�&�.9 �g��'���T��̅��틇jH	0}vx��>�YFꗢ$7���yf&�Y= 4�I�X�H�Ӝ�#�����]�h��xJ$����m��lҵؖ)Ӑ��3�J*
��g�Kޏ�,~rA@�tZU��`�;����B[�d8D1��0���䊏�k���G�˨[ (�wx�¤�ͪ�֗�M]F9�������HT��q��@"�p](�Q�k.%0����.�[���&JA�7ȱ�a�@ɨ�v޴�ߋ�ۛ^v[�VJ@�H\�m�QH�Lzߋ%=���
\@}���n�.6,���m(��b0�O�R�ni:<\�H��T^m6�r��x&��O��q8s��N��*c�C�z� amR(��T���Lװ��>؇�����'��}��'�IL���!�z:rYёXmR�_�ṿ)4��E�
�YU�4�>�����N�Q��W��`hA�`�mh!<9�_-�#3��ƘS�jEq�Q����@i�A�bI4^����?���O���ZR�%�w"��qV��yN��!Y��3�������ы��j=%D�6b1��]��URB{�7�u�V�(y�(=��t�
�!%�u�lN�.�W,7u3p�� dD�a��9S}�/���x�ܰ���*��̹n��}!6U�j��_w�*��Zu�1��-�t����sU*�]�*ӯ����� T�d@X�ܬ���hC���J� h6�|tQ�;�A�@��<y2�3*������1,��E˺�ˈ_��CԝG�l��Tܛ��Kr�����)7�$x�e�:pc�����W��:Z��?kX����\�Q�f��DOب��l.k���4�vp�s2p�4#v�g>���4Ҿ��|��8hp��ڎDa�31�R�)��C2����q���$Y�6�\Gjw�})�W���"!���܎y!Τ�"yg�y`���"��}NM����̪S�Rk�J
QcQ���z�_�p" q���lx4���oM٢ކeb o��x��{�y�e�e��Ehd��;xi,����z�̜�~��͙��)��É`q���=No�{�}Ӧ����AF���������AY�Ea"�fy�z�0qv��s���V'��f��I̹�pG�� �\T��$��-q ��WT^;�3'���Uz!��>3եC�B � �3��L��*�{+���/�����^�M9EF�]�[�`f��C�).��/s�NuJ󎃕�L�M󇲥�M\l�UTRU�6�擺�G�CX1�%���߉�϶z�g�o�<=�����kO��d�B R���&��'�O����ǈ��3[���er"��@�풷=#��՟���CXJ#�> �x"+-��R'�N��R�uz�}ǨfC���g(�C��!CՂ�+�;�C�>����Z^1j�	�iu*-~�$��f�y8����|�w���zA�RH.�R�����1�̛ �fLY8��DWˣc�N�	��EZ_�0�\�y�}-<A��Oړ�bM�W͏��s����{�(Y�ɰ���f�=/5s2���>
���ݺի��U4%g�:	&�	���ءB@}�xO&�s6�Yi���i����Eh
 �	��ƺք�F0����&6ǝ�F�
�ԉ.wK4m�:m����u���CtX�I}iE�r|��,Z�:��"Cʧ|�0�w����"�kTjS]��K݃j����)�}>�������.nF��3�l�18�k��:y��I�w�%����΂��vYhO�ޢm�VX����6�'<<]��N��$@uf6~/���h�͂����G�dt�_[��WA��ܭ�y�8c��w�R�{;��{g7R\�v��vZ�	X]���l�[M�1��0��,�;h�/}�8f��,��a�́��	�e�R���<�R��_z֠����Ξg���UJ=�5(}����)5��m-C�B:���"��C0n��j���x6={Gys��%��͌O���OBt8���nҹ�a�
����#��c�ˣXTz��������YF�W�0��H�Υ�p��(��5�8ֺj�c���K�T�E�z��\+ҧ>Gyv�l�y��,�31�s2@ǧ3�1�#������Ay�d+��%���RP�s�i�הܟi�O�п��ri��m幈X0�r��R�ybE��>�3�B��'�'s�>��7��J|l�R$�#���6�8O6��/�J���\��(IixP�L�A��Y���N�ӎhF*	_�
�I/&����;���z.N�>��F�D��Է$~L��-j"�v�A���?�V�Pӽ���7r��Ң�gl�q+����>�҉���!Bo����mc�jX������M_���9x�j "�q�52�9&:�(5:hv�	Z��|�^lS�Rb/��*����z�y�%R�L���C��`�?�l�:Rw��0%\��!��{,����j�F&.Yؐ���hQCδ<��xZ�xz�:(��+��<ٞ�(i���M�y�}Mύέ1���������Tq��{���:�[W�ƮW���v�#y�]`F��_V��Ĝ�I}�f����C�*�]�/���۷:Br�_`d#�e��j��ְ�U`D��{z̤�1�z�/�J�A�␜�|(�b1�?�8�j�݆C#d��	��>�˭�X�H`�٪ǘ�����O����|������ZxTx؞&{>�pv-��s�<��\�U�iX���S�o�T�iwG&!+*ʆ��c�2��C�E���l�	�%�WZ�4�t�R��ڞEU,I�3�R�����;�f:<M'�