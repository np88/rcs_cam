XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��{U?��{��%�O��\�X�����*j0�~�?nߢ���Ov�Ξ��czR5wR��o4��V�	C(�[��a���`z {��Dq{;�/�.-4]lL��Injpkr��Xn���lмJ	��G|�aV��3�Ͻ��WdX�G��RCx�n���M��s�FK�n�� �G�u��Z�?�w��E����է�f��n�u�� *|�ë1J|���7 ����9
���Xօ��:�xH�����
HYbZzS�:��h���X�͎+���מjX�ژ8$����jk����Ǥ�O	���'��D�ľ�"���T���|�Mi
��$�ITǛ���eg�j���}��}���5M]��|$�P�s�2���� s���S�o���_�,�}��岮��A��᯺ruPݪ�t����Yz�N�n���D��= �1� ��^vkbP�����k��fɮ�E�0+�{�	mS��n ����� ���}Q�8S���G?�5~2ٌ�&�O+�_lW�IG�FR�n��	� '!0u����k�� \�����LT7f^��8K�': [�7W���϶E�5����Y����号9a8��5 4� ;��ў����_�(���]i�K�Hϛj
7��ى�L u�q�p*����<?F��I@>v��;0!�h(�UiK���y{`�f��N�0���Y�YQ'���������3�nݤ�g���I����/�yq�fk}�#|XlxVHYEB    2577     a70�a�Ә�-���8~7b�ҙ'��R�J'�h�DE���ɋK�	xl���!�㈒%�D��9�?��� o��F�S"K6G>��n�x�Q�<SԠ�S`�m$��N����1�2T7Pӈ4CY���p��bU
eb����B���	B��/��e�=�#� Ѐ�>f��o/*�0
4�|�ʁ�Ԑ�59��!�y �{ԡcNa�	�S��B�z^��A&sϬ<����K��#7x�mH����d��A�g+�������IIi	��	mB��43��ϱ:���(y~1�k(+O��C��Q!�)�s�Ia?O7�͜$Pko_��j�=&~0��N6�y�8�T.Go��`�<���S���f��&r�'pf�4P��F��_|�Ƹ�����|�� ��QgtV�fV����-���.�:�a.����u�Dt/��;GT���\'h��^�&���ٯb/��� .��)�*7Y,��+>x�P�{�d�4�m���X&�[^(3�l�X�j�\4�J��������m ��ES^< ov�<���0����!3�r��^�=�M�r�%�ǘ��_�<��F%����`�\��S��/��f��%;��"�^�
DA�z���-��kp0?�ܢ���đ��c�N�����'��]�����(ͷK�L ��Ɂ,��Pӝ�$����Z^8�&Z�т^m�2�Q����6T�;>$$o;}R;�>������;�낔d�<��Sd}=���������*���!-e���UH}�h��#f�&���F�O��o��A���	�Q�f��;�Ʋ&ّŇ��"=~�|��UV{��!wE��8�Y�>{m���KHtO�b�3�,�
��,h/�����y���N˰e�����G���lGV�;f��_+��f�2 8`?�:j�["d��7�%�MP����O7�{��;b���J��\�L����AqѦ<�5�-�P��NP3F��L�$��p�L̽�d�#o�5�[�o�&�s����43&P?6r�c���7����*p5F���u��YO=�_`��X�)9S(���	�.�7y�_4!u!O[]�;� mֻ>���XB�C9��}/dm����Iԝ���j9��\��B(s�W��D�S���6W��*��,��n�WZ���P�Z[�1��j,ە�$�9ƶ�Eqe3wb�]�g�y7��H.+�<�R���{�0(����vAʼ����i�:&��AV�������0�:�+$d:��.��M�5�~�]r��U����7X��P�V�ֆM��/�q@��AEG���Lr:_��#�,p��������d�Xctc$P�wȻ#�5)W��a�����o`D�z>�3_a~�赚�w�5i���d��Ի����������\���'�)�����B�xλV���8z���'n�f��8z���j4G1`.�!(�\n�"ʹ�}��]$]ڡq
ZE�0�Y+���6�yaťY������٭�l(G��oq����#�@zm�P0�Ui��-��wJ��H0�ղ����	�H��s0�ĎTQ|��A�[�R}���˰�<��#,�8q�G;�"�.�3�'�H/U��pqIW
z��wb��F���P���)}��\[�)��:��ݩ�C̀��g	�Uv��n��R��dh`�����>��]��0i0��R���L���
�M5����'���V���@E���_���K�V�[�"�N ����O�Oc�q��)� ���Đ��|
(�[�Քޗ��v��C�5���-��}�:�RbAP2��s�"cu���5�d�b�h$��X7@o�K�%6s0,P֚(z�'���B̻��v�[P�aq�wq�HsI랶2 ���:H����; NVR�
�@���.M-x�]/��C�Ɛ��4�����iw�NRa�+�1Z��e:4W%��a�������u�o9<�~�v(���e�8��pAH���	C�����d�\�{m}O���&�p�9��&�3����.�;#@�ԁ��6�E��xƭ(��D���@����P~�ZX�<Yo��->��4M�F�<�(K��B4�V��������^J!NT�C$n�lpP(E�D\������J)�<{U�
�#��4��*#�I]�\��!cEg�Zǌ����jq "�w 6Q�5V�#vo|��6���^�����AF�V�<���4���=z'9'FU+z��Ç�����$ �$Y���
��U�K�^Ķ�ۇI�lHm�J��t�_O��;���	X�_ ���.�yI~�	�D7��khp�A~�mV��m�^�!�U�+{� _|�����z�`���P0��T���qL�hH/���q�Xbq�$��5���9 ���`�!h��EW<�.����f�s��e6�N���6B���<.���`l�ؒ!��QE�
����I�Z��z�z����Z8�J��ض���ͤ��h��zR�W��+T�Hh͙ds���cD��I����!��d
e�4�ٸ4"	�Z�ך�
�'���mj��Y5?F@E�R[3	|W�&9*��V�D�-����T8�a���J���V���PX�ʄ�ݴ����
�I��E���؁@