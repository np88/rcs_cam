XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����Ui�֢K����*�\_y��=N<���)R�wn��Ü1��pz�N3��f��%m��[rb���[�s�3d���	z�^�nm�ŤAk�M�FHm9ܺ�#>�+��:�/2�ζy��ξ�N�Ei�t��&�
���V_c����(�"�Now�<���ߜX]i=��L�C�EY�#���.���x��E
f:*zv�z�Z�JGq�V)�t۟�$X{o�2�|"��Y��7.���}��}0� oY�����_+%/�!�D#�z�N'G�˖e0"�,�lW'뛶�4��u���cV�� k���F��M݀����<���n�aM�8��פ��}�a�e���"j�ȓ!J�Ԣ��8�|,u��;�_e+р ȡ���.�U	�{δ��' xDh��z�����9�pA�/�Ÿ�����ٞ�(h+U��uTT�(�Ҳ���ZT)�CB��ۊq���G���V�v����7ށ���0�e?ĭ��?Q�@�&�ʬ8lGIpPh_��V�!��q�y�����3/�M��3�!�!b���@R�Bd)��v.c�ۑ��J(;EḰ#�u>v�r*�V��Ӑ,�58��f-UQc��I�@t 16����3VO9�"�����7f_�nY{8#wp|�G���Ÿw�FZ~�M4[��ԇ�{���	�2}��e�y�H��Ӆ��{[��¶�F-�@�pk@�im$Ek*�(�Wbb#?�\~n�0�6@E�{g��򅵤+�3#v��},�	�%]��#:XlxVHYEB    fa00    1790<�|mIi!�8㉆4��u�IR���m�5�"�x܉��b� ��������Κ����Ң�^i*�_��?� �fD��<y�B�� ����tS��vhB�/��Ͼ��(p�2���x)�����bЯ��Wt� ��fͼ�aL��xU>���N�o�I�+��b�8'��DPN%X���2G{Vb/Ԃg��Ś�CS��{uu<|�8,�^�T�"�UJ4�i����������קF
G`�3+�%���+*��CX;x�d�ٕȤ�#P2�3�S}��;e|k�>�5���Xū�H Ƴ(j��G����Y��%�MR�n!�{��DE�s8��l�̞T��ՙ�_�/<�q��F.����3�g��O��j�"��cm�u��z��-5���8=�!8N�9��n�9]�8���Ce�Ȅ�'�L�1v��ἧ�Y�����3zg�Sc����M=snh�#g�'�/��F�+�/X�nY�1ݓfg4�RL��`� h�#@W}U�<p�6�Јuf��"}8�2`��a�K��/ִ;M/}��M�����B���8})߫"i�Eb���I2V	�y��N0�C���#�Է��m�.?��Ԙ��축qF?-�oi3��I^=d���2�IK��^_=؏?"x��O%��1�Q�y3�pE��Ә��;�u6��L��S�!�BM��Qym�C�s�0p���,��e������T)�����W�%�P�n*߫mt��1�/�˿Qz/��	�OPʜ����<&롼���2Kvo��!_q-3�tfU����u:D3�2;8f���>H�V�h���U�E�L�%�a��c?i�q�v~��U����~L6Gk�Ĥ��%b{�n�S2�O�l:�*d�]-h���D�c؈�ܐ�I�-M)a'>9P�����d�A�k�x���ʈP���'aMs~���x�J�ۺ�����6�j`��"�NPf��]_s��}6;��9�<��?�X��W�	G�����+>A����m-��e-�ar���n����HW��y�S=l���dnP�w~>
��x��	�N4�XX���5
�u�a�2�����Pv���j#B�RG��GX{*A�E��nU��-�n!4���mG���A���-����F�6O�H�=i�̟?��L���� v"�D%��`�P�_u|����))hȷ��P�ž�h����'	R�ח���
Ӧ�YA�
Z�_Y)@Y6IpB��>[O��o���W�q&��@���������;�#w�����d�n����<���i�]����Qզz-t������{C�8O7h�"er� �3+�����fx���;��X��ᨚ�Bl2W�{�H0K'BRF
ً�7H��=
����c׀�q�,D�����i֖�{'ђ_ �!�}���r���2$9�X��L���7�.�Y�k��+����?��(e��h�yeD4��޻����o=B�hvik�_��Zr|���M�ac���
+jۭߵ�9�H~�B�r���R	w��8u�hY���^y��Sb�;O�|�,���?����o7E�Q���%k��QjNЗ1�X�t����2��������7yY�8��%�E8w��h�N��z� � ���B�!>���P ;j.β�Wp����@�F�#p*/�\�X�Wݖ�}��JRe��=��<��k�)�'�}<��Ȟ�ڂj/gq٤baP׿��+���.�1�9��M<�({���H�5i ;�-L�o�����w�^��oϰ\Q
����������6�gs��E��K�YI������sJ�F{݄������G��+�q�/M�;���m���SP�9�h���ԓ"|�ȟ�V�����1�$'�f�ȥ�ߘ��uj��V�$����^[�U�2O�9#�X��=�z�I��6�QOf^D�X$�*��^uZ#�tu�H�%Mɨ:?��&�.��.���NW^cߞ�������T���b�k�)��p+�Y{�ñ��"�?����џ�9Vt�k����LLn���K�*�A��VgFk��xG�j˟Q��ryvuI΄��c��=��;<s|�UK��p�t����Z�a��W&��QPu��u�߫�G��ax������'��
<���4�hA)�S��*�I�J�܍ـ'(����A�<�5պ�۳R~�Uf�0�2����݆�u<�:��q��P���QX*�z�2���4�w�L�T�طQ�S��|Y�[:v#9>��jJ@����/�q�m���yq!#�l�w�e�U��ܵ6����:�q���VĠ�9�E�LE��֙�FY&�O��E��W�m 5@/A��p々��R�D�n�ԁ�V�Ty����o#��JE<�AJz~f*���]�N2�/��؂G�N�,�7� �r��k����l&(J��s��L�O=C�|Q��)I	b���Ɲ��Tq^�sZ��|��}-�㶘x�[��_�.|�%yJÄ�҄��	 E5%�$�HCs�f��"X����eP*f��.�?X���w�͆9E�.�)�l)�v����t�o�4�7��2 8T����z�C�Jhy f�׀���<�0� ݷw���dW+��َߘ�H���y�/0��9n2��~l�œj
= �Y�3#Ȗ�P�0�[��U�=�_>��25�2�7r��	A>ܕ먪Sz

s�N	+�M�%��=��ku��������R�%P�~�I�1��,��s����Wך��F��O�TU$)a�M�)Ic��p������qp��v{U'E�]M���?s\��HE��Td)�]$ �xX�b�,��~�
��[>kej�0�X/e�p@�!�h����bZ�X4K��6�}z�#�ه�r+;�Q�vÐ���ƥ�}WM�lj6���SЈOԒ��hྼ��"��k������XY޵M��!Я�V`!q1~�>=e7���1�<ҝ��*\8�>(��Ա��Ê��C�q*��,i�JY�a2;eED,}�Z!��t��& f��|b�d�є��eh#�]���f�q�H�J����2u������!���Nl��O�;��+Q4*B䋱��{P?T�	��&|c�V�6�Dޫ�����u�"H��*a��I������������@��r+��k���r�x|����^������J}D�� �j�K����v���Y����tAh��V�d�s�)k<��sİj�����k�+�Ƙ�6��?bnɍFt�Q/�m�R��-����_�s_�[�l�a�"U8B|�=RrPo���zό�6�fFCv��T�8�w���Zk﷓o���:z{ F��*�#}h��M6��^�(ҷ�4A�R{�\�e#'����t�x��I��
�{�Y�Ӡ�&��-#�PX�%�Ɓ���ѸN�l`
ѹ���[��?񟿼^�5ƪgy������,���
*�>���aS"5�p� =�r1�[�m�(2(�V=�{��������R�h�f���a��r��0�Jv��f�N��Z�O�$?�×f��Vqq���X7�ȱ����G��B�}gN
��K{B���B)�,`��8��]�t�n�<�˸�
P�,�@x��md%4�0i�����sb��4��*TԻ����mt�1��H�F�򪊐,5�O���h����`�h�O2e�x28�����PL5-���G�Vc���F�˕�Z"�R�i������� s��N1���{���� �s��xAx��~� ��"��c��s�ȹ��Q)�z���c���Eo�O�,DZ<�ϛB/]O�~��0��l��S`{��Y#K�B�"�@�|7ʤtW �}�.w�_�s����aG��3�*i���
��U��mڱ	ĚT�!h��7��5���'���eS:�O�x�!{I���dTq�;Ȝ�����"��c!?�
\(��
��r�����-�Mq
Q˸�f<��l{�C�Ǩ\(�fٞ+?*��r$NQ�"����c�s96"�5��q">��8�v'���}.b=5$�-�	����҉�'I�Wc��45�RE�Q�����&5�0��G�p����9��v�d��R�
ry�pD�,�g���]�Vy4o��z�@�x�!�ҕ��W��R��2��ɡ�:�e%=3�꼙��E���n$���7%�_9�=���`M*0�0bE��$�T���3�x}-�Ʒ����RR߷���<�ζ�uX[�[
 -�ӃF
���4���e#��K����#T��Pi.'-V���᯳ﵹL󬓹:�9T��~'�g_o�Quz[k�hFqfNؖGA�ⲘY�v_8e㐛��nش>zn3_W6��s�� W�,�$/'��t�@{L\L���8����� .3�u7�� K��!���d*E�w��(g*����umO)��SL ������%e>��!�<�6@�L�Z��
�C�X�g&94�[��*;� ||�Gȳ!�䵆�����[}�U5�_G��'���]C��E��_�Ҋ�[d7��M����雾�]�*�h��d�m5�����)v7���I{Q���y�jR��.]-	�o�Y�}�P�<9pi
k�;���|���l1u�W�d�R?Ƭ��'F���ޢq+a��G�����n��d����8ę�=��~va�Ek�y u���6k�t&\����qx��jL�>?��M��\�n�;���kw��p¶���Ư���::q�_{���v
����'>KD�$:X����4@�a�@�U�訤x\��`����]�/��=�x@p�ʜu�V�n�"�n̶+�����&�m��$�o�2!
���u��b��FiYZu���TK��$�!#<��R3�\,u����#����pۃ�C�!�\aE��iah�l�9����.=�wpʲ�q�u��m�㈤k�� �4
��6���ڼ�D�2�Yq�̺ǩ��3oi���2MQ��J�A�����Tt���4ۡ�#ā���j竸�:f��N@����ٖ/E���{�T���8�V�X�o뭩�����ڵ���(q����X�_��'Rn��y�D}��j��/�Yc���Z猾nI�
�9�I21@�DY@���a�k\a�5�iv�i��P�w�0�M"RH{��諊б<N`�g��VkO*YP�'����5x�bO8;yucS�a�
t�ɉ�\:V�fm�R�[������'-�d'j����<q!��ItU ��Z����+�� �����茽0�ID������~bq�8\���Z
v��moӕ����΀�w��D�`��'��� �T���9%�u�p�C�x�^��O��#��磳�J%0�.[���a�%�� ��)�JԄI/ҀJ7��e��C��^R�������M�
�c��X)�����G��PȦԄ�,�;c� �O`���F{�0�����_7q�#S�	%�j�?��W��ZBC���-�k���ͭ��x���AS���\ή@��!���������@�Nq� �Y���.�M.�m	�8A�G�	����,���9|.L�BR!]�@�03F�x{�3�~$r��5��2�[��0��1�	X�E|lѣ���"&ޅ�*���^X���r�L��'*Bmh�-��&�<ۉXX̤7�2!T�u��*�� &?�s�o���..] w�s��c܉
��DN~��ɓ��;$&�A�0E8k���e��(?��g�X'�.���wd�ͺ�\��ah�M$�s���RLrV�f�0��z�G#a;�3���Q��@ ��3�#��ϭ�\��>L���_#����4�r��h�d[�[����ٱK��bzJ��Wӎ�Q��	�����*\�1��6�.,[�At"����Ԥ�-CgDا�F/"�������>��-piLNx�F���&
a^4������gʭU�r���BQ��XlxVHYEB    fa00     5d0�IQ|���,���~��$����Yٰ;�^�ed�7OՒ��q)V�.�0O��o�P�u���[C�;v�� �07�
��7dN:��R�A�/�2Φ���-���ʮ�Xy��)Ě�������jW�8��jCw�0���a8?�R�h�6%&}c��b�l�n����&5u-p�<T�}�C��ސ_e�f�.Ji�I���x��'� �2wM�1���N�T�����V��Ǽc_�RQ��<L=��`�]`�c�+(b��d��	�Ce<���6�ޛ5f���C�~��G�a��C�p��n������9�8��R�Y�~�p��OɈA�a�bnc�P�oB�/.��.���C�j���3<��� �Ѳ!`�:�6�J��;�Ѯq����p(��eT�瓛M�\GAnͣ��P�[�~���^�7�5��Ga������V�>U9(HF�m�	�&1��I6��)F%"8�����W�x��>@ё|���e��o:��߻��>c(�����lAp�1M'8U��}ئϪ�-��ut�폃ܗ��lc�/�g�uu��C�>s�[֠*��Խ_���]*���|ULi�3xO�L!H�_�v�r�2Y��柦7�<M�kQ�b�9��oG4���R�g7q���B�-KS�%�>��f���yr�	�'����A�r�+��$��tN��%�cY%"�gI�n�i�[?�)�R������wݓ�+��v֟�(;��Af�Πie1}X�~v��{�8_q���]h5�͌?ƽ��0n�Y{a�ID�
�zQ9l���w�Zޘ���W�<(F޶��8�nE��T�hM�K�2��ko��B=3�1�CŲ �Q��"<�˃J�JLT��S���䶳6���C�ѮH��E��.�*Emc;�A�~u@��V�E�u�tU��X5�ډ.�R�[� ������� �#Z�q��_�f�UX�Q�$�s���]Y:Nyt�$���4��
rL��߲+��1�̵��?�ƻ�ř�\��k���f1�\���/��<+jԭZ����g��a[)ݩ�d�T"�Nm�A�I�/�";Ut������	t��\�E����K�a�?Z�o��B�3%n��x�R-f7��YC�>�n�\W\ڦ$7�9 �^ !�;Ax�f�~�۶�e���˼Y: Wᆿ�y-���Ԉ̰m�d݊AB�ہ��H���C����m*�8<�W��=&u,wb�:�,��Q���|���G}���1�!9gҧ <�Ԋ��ꍙ�����B�/©N�k19��Ղ�,9�@��K�h���fK��>����!�˄?�9��M��_`����x���P"FN󂙴R1�j�6��K�*�&��q�B�X�2LLT���40ʴ�ԇu!�R������6��Ue�A� e9�'Bf7������c�!A�ȓV~�"jr(?��]�(jt�xVoֱw��O�8vBIRbO���XlxVHYEB    fa00     640�zM���.;JN�&;�S��&��+�K1<p Vx=�@]�0PѾ^j����HN��|�J@[u�
Q&ѩ�!=�]:\������g=��*��P:���Bk�Qr��p��a��_X]{p��\�l�hIkT�ɰқ��$ e[1r�C�^Ԍ')�F���R����yR|�g}������r$k���X)j57/'�RQ�������?RXw��#�>�F?�I�G�*��-��F%Ez`�|�l� zu��]�큛$_���YG���F�+�����;���{]R����W��3�D#�W�I���be�g��C��)����
���d�_�6�CG2n?;�I�t/
�Q�f��� ���N�E�.����i?��a�tΡ Έ�%{%�{;�c�y-����K�X�m�{de�#���D6Q�@�f��͑t~5p܃����ȧ�U�>���g�ܡ�.Xh� D�\��}����=� ��>T�� }BE�؃���P���C�\�l}Ꮈ>��ѕ��F�z��tnL�@7
�A�onvэ~)��ޱٹΗ�찡P,b�ϸ���0Y�ĽQ�����8����.�<H��L�=�b���1r3��f!�{Dړř�,+Y��;#<�oɖ�V00��j�'8c�F��!�>êq������r��#��L�C�)ȫ�= ���a�(N
˗6i�E�b�k��(o(�`� t!��_j����FU�m� ���/C¤\���ީ ��	����4��s�Yr%�a�_r��ƢGTe'7_�(�>EO�}��5�x���ȇ����wK[VEkx�0���,+��C��B���у-�>HH�/T\Ö��eG�-���g�i����8��&/�5�dϝCDiAMQbp�5"O%��ڗ��ez�G�ѐ�#2ތ�*���F��ܗ� !A3����9d;H�ľ,�����ʋ�9��O1���^��L�^�=��Z�o�̩^f�!����k��l�z���G�/B/�`��k}8�AG�Q{Ӗ��t=�T� �ý-0'Kyx��n��Lj�x�o;8Y�����pB6�K9@<�1h�	s��1	��yF/�1�C�C.J��C��'MCL�����F��F�1����*sUy����8�{ �9�Z�d�����k8C�� ܌��ƪ�׺�MVP�fdF�G3ڣD?�O��H��H�����*i�AÝ'�S�V�XO����\�!Q�t����6�*Z�)��PR��S�A��-��4�Ǆ1�ae���>!O+���io�c�j/;6�����N���~�F;V������)q��H4;��n����{� �����F�2玊9�A�^�� ��EW�����J�zk��?
/�j$��5(~�N�Y�.٧��T���w�%��Ae��W�ѥ[��K}�b֞mlO=�s����BW�D*v�����
D���RT� D�_����u�"�i����Tvϰ��ۋE+r����k�]s[�IFI؝�4��P�&�n^	��uM�I�z:�W��O�R�Y�����+DOm������A<L�D~�Pt:�x�G�@auJXlxVHYEB    fa00     5c0j-b�U���=�ÏUn���-��$��9Ƀ��W�/��l��b��LN�յ@��x`0ݧ-�{�
)[���k	��ܬ���Q�Z�z
G��Lg����h	���R��D!��������?�����1ي�ɭ-V� ��yek�6O#�B��	=,��]~��!;�o͚��I���f��O�Wo.+]i�XȞ�c,�Nh�4���"�v8���n��dl9�Ά�"�WT`�U2%�θ_��a�2m�>�wV ������qo�ic���e��(�N��)�@���9���̍A��<��}"Y��b�l'���|O�����.�SN���1��a��n� #�3�w�C�5��?[�q_����g��`	W{�ې8�3�b=$#B��e�'/hr�����ID��J����U��o��}�}�lrx�e�&-4��]�UR�^���J��r<S��A�,s�l�x^���W�Ha�	�S���]u��]֋������.UJR��olp�i>)���h��n�">>�#HW�D���)SƓ|_�	�R�a����@}����∲�ܲ���w�3�����|&����G`�o;�af���/�:������ g�D��'`�;�ꆾf�e==�V3�U��� �x@'�G�ދ�����4ۡ-�!��U�R^�������?L�f��#HY�V�U@ O�)s�$���1=�Lv�T������$���^)�����`/�3�þ�A��>�-��p}��g�&O��;�[�U�j�a���(�*:��N����?OQ�Zz�i	v(��BV�jǱ��^�̨�0yAk�+E��hL: pE���������� �*�������*Y�1y��˾5�Ix̫U�:\�g�ͥd�q�9 T�� P���IF��;��*����W"�β�OtR���N��ֈ�2�쪑���Y|��UAy�e?�%����)Ȇ��;���em��@yʿ
Lz�i��1p89��^<Ȭ�=K�a�)C&�l
���Ki��r���Ms;��U�**���9���{���dYۉ P
@;|/��'�z���2����Roc3*���S*���-Jz�(��c�i{��� Z �Gf.'�D	t4y�3̘���Ci��_�<5ק/�m�#��G쯕�){����\�h /cpp�,I�ɍ|B�>@�L�f��$�<@��lY�-�#LfV������TA��?��D��fGCZ	�i��ݯ�q������)�����hT#ʘ~�_��K���ٿ4�ܾ���f���U�t猙�i����5�������>86q��Ϯ
0�G�WkHT��snS ڋaO�"���׿M:����	l�}����q}C	e<	Y��Trr�-���E�ß�{=�'.!Z�?P�`�rU�
�Q��G����P:����ɠo1�MXlxVHYEB    d347     a90u�o�U�J��[�L��I?�vRs�_��E����!�*��	��x�!h��?��f��hbj���Q��]Q�`��0�B?W7���c���U�y�ʩ�.ܺZ�s3�x�}F�U�_u|o�|Jz�������T"}��Z r�����?pO7q���<)y|Μ��%ئ���h��z��IE����f��iR��g�FP�ɥvGV*LH(V�*	��L���]���6��`���q�]W�$��"�]{�1g�I���*]q`� mnHy �7 ?H;������KK�m]�3g��۔%M���(�-��K�,�U{$�g�jk(@y�&�H�d��1p��ir��ۏ̀ɝ���|����W������y��!D6���V_R�0�>!n�u�e���wY�v�!��A��9��M���,������� h!�3�ء%���"v�����e4J>��KG�Ն���e�/�]�"���z��su�s@�-��<��=��x����i6��Ǧ[h6��ņ�U5\���t�.�'�߃Y2g�a�$���gg}����~V��/O��te}��][+�6�(�e^�#����-nRN�"�!�2Ϧz�f�A�io*R�h�����uj�$��C	���Q��hT�Zz����P��K������u��{x�mc�ٍa�8��=Q4���膨4_���Aa�O_�#��4o���0u�.P=]�����XFib�V���Qu��nx%T�1�ăj��1��iѧ��'p��y���9_+�2���oG�xo��RD*�~��I3�&�W���M�8ϮD�B|W7o{���>jN���z��V�g��������c-�ݖ��0���ֻ1��$�7�k�ɺt�?o��cNJt�������D���q�EN6k�`$��"���Ko�����6��o|�@���uZ{�m(+4&�n�ph��w���y�$����"L��e>o��}1`�-�����R��G��!XV��n��B�ؾ�� �-�>��dF�E�:�Hj��Ǒ���k���i>�� ��5�Y��?$w1��@���:��PifV���T[	GA<d�����k����j�M��:�1cW1?�J����FV� w��g��mpp�����{�_�� �jҌ�����7S���H.T*�uZ���V%L���).f���|E��m]>Z�o�dxn�%�@��(ǫ���# 9u:e,��8!|P?��ɻy�(�錕���ר̅�$d�R�6�|4F�ze��lt�I�ȭ��q�Sf��;�O�=�A�@�Tt��,$>�TX�U�%r�/�s#bݝw4Ƣr0����&��1p�~��]1���2/�
�'���֫~� ��0���7~�9J�Kw�����U�)��U��������$��w8��Jz#�^U~��z�hb	 �N�o�VR�z�\�|2����|)@fۉ��P���r�S��ń-�T~iթbs�U�V!�h�Q��|n^���f������v@���(���u��m���E�c��������E#����7�� �ٲ��De~$��9�6l|F<�P�*Ѽ�iy5�����hp��Ah+��g[��G��=×a�s�[�c\��`�fs�a��nP���8d�W�*��I�9M>'���F'��o���8�m#���G��j�W�i�x(��m_�R������$6�B��\4�*�q�k�a��3���ζ���ƞ<�╥�h�G�_T���駴��4�:���g�]�EI��o�rn��Ƅ�(�p(�.�G�Ë������C:���2.����t������y�����S,ЂHL����_�y��y�J�F��<�8��q�o�m�(˖]Zr�Vz�iw�����*�ךD������|f�QL��Qd8��?��Yhm�Em��[r�,�E�`V���O���y�AB�d"���>���Ӎ/��6��d0���f�n�;�?6��]鈋��t"��Y��3 B,�w<d���/���v(>s���}ȫ�_�fC\f`�2wW �D��  ���������C_�j����2&�7V2Ez�Zgc�Q��,�`Q��g+g �ubpP�~���ͥ/9cd��Y��QtE�F7Ⴊ+�k��������#z�1���L/��X��\��	�tW� ��
��rui� TO�_t�:5��;����53�Q�90KժH��J �cT��H?Y�;>;p��n�ee�M	��*���U��A��tL�&��{�4��6;��,nv�&cx��~�]~D5
��g����:��dS��ڝ��a�WƯ�h"�.SN��Wpj�ۇ��f�^��8�#�!V�x�{���HL�������ȽNS�j��%�����YT~Q���H���USK����3;Q8�8���:�j�����!W�;n�;X�ǹ�p����Q2�z�o\��=H?��9�`���Q��G�D?��fD��q�{���\h��T�ٔ.n��\��6gW�?~�y���i70�S	�2!l�q6
�(ޝ�he���;�46�X�"�����~��4��!�xY�����:j����:���h��5<��n2�r�ۡQ����`qvo�+<�?<�ޟ