XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����
�Ք���-�A�ff�" ��l�
���/�����L��_�Q�TZ�>��@p�jej6�AX{r;W����+g�V#Vof�}�^�A��e5��$�(�fr
�������`���?A��s��2�%��5|�a-fbK��`ojᖫ��JѠ�0Yj@u�T����N�y's�P>qb�_fsy�" �0s�z#=�,�2�����3� ����޶Z��r��{5���m�풹=���ュ�}�J	B�Uh/�Ȯ,�X��;ڇ��pZ�V�#���^�.�'�q�>pC*���j���d�;�R�3lm~{�1��6<l����
��:�U�6�3แ��{bO F2b9�x"H8@����E��vim���C�`Vq�T��}��!���a�h�+����s�U�m�*��a�h Q:v��LX_���,�.MC)8H���>s�=P���6��#�G9Ò�J�a���=	�rE/� �+2'��UP��E���֤��#rQ���z�.��-?.1�
��͟\H�JR1�fd�]xr�[� $�A�(���ZV	��Λ�1��&��-����m%��z��@�b��]�̖$3�1�;����yw�(a'�#%7�@�a5Uf��8Oi	ԙ3�uo x|����ey���r���������Ln$d�\r��� k༬��İ�#�Y���`X�c���i�8�iH+F���<�?3O��?F���ٗY,�K��*��For��j�C�s��e_�)6����z���Y�a�XlxVHYEB    2f9f     c60=<plh�~	�(
�W�<	8b#���r���c2g��� ��QX7�
h���@@+B��,���=���� #���.��(����$}x&�,�Xy5�t��S*Y�a:Snڂz�9��"�C3��T:Q6��U4鼴^~����G�9Aݯ\<@;���|�~}� �r�� R٪�l���+=�*��c�ݕgBzm����*V�/R�2ÎZ�&z}D����8�:,5a�ϩ�
���Z�&�g��0:�)u,wg�?9�
܁����98͢�(�myU��EB�� �Y�z=�_N���W�H������5޻���[Z͓Bీ���݉N��F��I=E���;�ص��<�=��6Ζd��z����+��l���r�:�I"��'�ˊ�L�:��{284��s��u@d��
�P�(;�-^ԛ�hj�guFƔp��,RS>AqP�*N֑��	O�kM���ZZ=�]-�~(y< �o��m��_��=I�<�ڮTꞮn��)W����o��LHy��v3�lk�(���}yﷃ��胲�����^��%`��䪛p�q[1'����uv"|Z#�P �X��Ĺ�=f�2��L��S����w��M2@R(����������\J�uh�GV)z݋×=�f�g���I а�b�����=Z��Yt�K���f���b�vmh�!P>3�מ�������{�@|O5�ȗ	S
'�뼟 ��K��m�Dnш��$Eٓ�I��6Qo{�P'Y��>
[��rB'�*����0��
E��:���� �k�qr��2�e�~���e�f���Z�������!��9����(O��
�Ih|oѱ��7��Tn���i��u�,#.��!=��2�M� f7/�/Ɂ$/G����NL���>��P���̽��0l���7�)��'혎��3jp|�-�o5�����a�ע��8�n��^%P������"��`�S'��oN!^$��Ϡ��-| O�;[*T��:F`��e��4��+�Flգ�?~18*��� �c2	拯��[�">)�ET�k*\AG�l[Bi���V��8���+{+h�oj��d(������6�`�M����� �H��૥}�w6] ]�ຼ8�Vn�Ϥ�
�0�D^�1@b����D�J�P��GJL�0�0�FXŉ�� ���
W`)�	���o�A,N�P���X � ��G�In��ϩ͔�X��g����^�+F%,���J�D�Ua�\̵XX|&��Ä�e�_���jI�m�Η1\%��m�>�8�߬���9Gr.�N��Lz���m�v���%d�[TVK1YF)A�F��&K>C�M�K�C_6'6!-Wp�Th��ÉK��B/���c�
b'���3�g���܋���w��/�����3M���۵PGv�~h�l�i��lfVJ��)�fڤ\����y�|���y�L�/�0 �
�w1���H��.��\|���VP<����>ř�d]���av�%��<̯4}��
Lо VA[g�G��vh�o���}��n�~�Y1����
|�l��2�H���2r��2���H5Ҳ�[��}z��?w�k�mR+��ȇi8��Ϳ��69Q�.$o���eB�����w����*d�A\��bI���8S�6��bܣs� �W�$���E�چY�hn�K�����S��RnNKHo�6��zŷq�貦hq�V�{q�eZ"�{�?��޺���x"[���.$�{Ads������Ck��/}n�w���7_M:îj_�6��)���g�q���ʌ�����ʌ1LD�l�=Ѣ~S��qI���̝��S.��P�@!�)uf ����;��*�2��1HY�:_����*K��O����_W`3ul�`M�Fl���a�O.��0h���JR{]r���v��N�\J$��=����h֚ń6�S�.Zl�D�Z��
�﷎HԼӜ���6�����/~��9j�O9ˌ+_k� OQk:V'z.K<�:�J�[O}���MWar���]/ѡ�V9�`�[�k�brov�EX�v�G� "��8y�"Cl>	�!Åy�U�Z����I�qv��\n��9�o���[fc���[EX�|xm"���r9�,I�b�c_;~�N������1�ҋT�=d���/.� �uR����;L��v�����'+ �I�m7ʐ�O���M�S�tZ�"D���f��~�m��%������f�d�����IL���Ѹؗ�4p<08��J�)#��F.�ˬ�"Ĩ��䓜��;�_l��L�s�
S��]A1H?uU��v�\�+"U�GE�C6a�V/�h��͒,f���r�Cހ�;�s��������?���1�M�!�$�_����=�����T���"��
/&FN��ߵ��y�G���� ������m8;�V? ��H��@�~x�����6}V~(�Go�s��!?�+�6p}Iz�/ m8��Z�
& \DᓋOn�]�|����LO��<Dh#�r����Q�����H|\�a$DTe�`�&�X~�A�,����5�Y\�G���B΁��$���?7q�����V�C7T|��P���0Jć@��B�cM9��ƪ���l{a�GH5��J�:`O�����_�mExςKE?��aF��C��ϐx�ʨ�<(��P�>Xk�k:mâ��K�w��?<��Ϝ�8��X}�I"
���k���(_�٪MB��F�*�~�}4[)5Re�ĄA���,�߮��)k0���U)�R9>f��-d��f%� Jt��+5��tZ
zC%���kpu�$�e)i���ډ����`�\8��f\�)�Z\�P���reF�6q�SȠ�tBb�� ��p�itT�s�:�'/���?]���z�	{�T!h,���N���\6���H=t5�\��D*X5?�[%��l�)}��VٞP[T�M�p�����~<����������5J�浊�T�%b|��SV�=�M⿾w��!��"���?�-|ښMm	 ����B�����[/���]&��;���k,:�ݹoyc?��=�����/���ܗ�x�8�fWtyR���B�Fyo��7�p���@�ke��s;�x��t����(^{�⎇