XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��V�wF 2A¬�䥹@"2[��J�����7�v� �	�i@#�P%��jV5��q
� ���oA���� �_.t���0���q@ⷖC�(�T�̎Rd��=Ta�;Q�8�����v-؏�1�0 �h���N�����Ý���?]�2yGi�E���~�3=�6�������;?j{pX���/T���ԫ�>�,��������������e��ba*�EO�Kb�޴�����x�.�����G%�@L8i�"tN�C���P�H��P�v�'��J�H��y�����m��Ԛmp�^�:g5�Y�>��Iy:��������h���TLOd�|k��d
��YK���+pē
��qb����Q�f뵑��)�Y�z��8�h�h����6nI�X�o7Emz�f��H�h!\���d�8���AS���<%�'�L�N�S�oA�D7hI?9>%�u<��h>0�Ju~ɞ4����O���z��A�iN���H��1�2���m~�����|�N�aJ"ʵ�v�h�\���n��=9�3K�s+�ł�L��|N�ٖϩļ�HK��#���R�\�g��a9 2�oҿ����	���kWw��5���/�)/���3.���x��p��Q1����5or�	 �N����/ϯ�>�6��%�R?�j7!PE�����@���3��٘�4_�E��ʮ��So���G�#�Nھ�z�>1 ������ՈU�.@�*�˧�|Dx-�jͬ>���XlxVHYEB    162c     850�DReAy�� �HR4%9_�T�~��$]I&,���d�>^A�"�q���,���y�2��f��;U6�@��c��X��^���R.�N���BD���e�!�{^�5x9}�l'c�6��3��|L��)Ӌ�x[I���=	�5�i	� ����&>��CtL�q��\��u��C��:�/j�W)\e�{�WxJv�+�Gȥ�f�&́6�U�ʖc�w�dӽ�n�@��8�R����P�KiHk�;�Q="�:�=�/�k�~xp��Ҭu�́/�^�2*��l�8���3G��#OS�_�23M����� Bd�NP`5E5�g#s�����v�Vn�,SIPV�ɇ���^� �pK���.�8O�����
�䮁�1�XK�����<��}��fgɣ��+Y��8L�}����oq��uv�a_�MK����svל�d�#��ˠ8�6-����`��_�v|�OfHh|�Д{=�����d/�H��<!a��E>Bt��n�#0%l��ٽ{u��
�й9�A��:��b��~�q���~[�bP�䰧�u�#��P2�#S��vzy����}�|܉:Hk�z�L`�/D������(
a�KBP�P�Bm���@����a�I��W�/s����o��j_�씆Wi��G�h}�Q�dRޒ±;X)c�|X
�s ���kL�G���o�<��H��[Y��إ��R�G�ิ3������Q��G��K�5�:����
j�g�ۮ�g2Ï���orK�X�18"�Bލ���N��d`��1�N�����w�4��>
r���/>S0|%uS�H��g�>��ĄZoY?�%���Q����D�C�׭�ϲڵ�s�1k-[�SJ��=ѩ*N�ʄn�8Y)�0z�a����PYq��n��d,�����~{����]>1a]��i�
�܆sTO�&b�K�s5h��s}aVt1��\_��%-��N��n�(A�a*�u��!�82R��j*��)��ۮ��L�B�z�xǹ� ��e�0���𜛭[�TĮ�kgfyW}��)s�Q�I�bY�y�5�8�ޛ�����8w�ȍ�QZ���`)��G�.�6:��F�J�c��8��fc��7�~C<��GF���/�kl�"+�s�kc#������s���UP ��9D�7����B�{��O�`��T���׬��3�
50ҋ��k��v������@Z>�eZO��-�� ]�3��%n�^�y�}ު����hFi�1e���?�j�)�ܓ֔:�
o4�Z����h�0^�1;1v��J}��P9g�>�4d3�$,_r�C	Ck;B�ˏ�v�;��-{V�M֒��JVo+kot��b��������志�o���O�=h�IU��:vA&�6���#�%��p��ی�芅�5��Lߥ@>6�q�ϥ`*��K�_s��`�up?w�\�4L�OƏV���E`y���I0��l@����ce��g�(�<�V�cF&���#�SF�Vnl9׺K��i����6��q�q��`����뫅pP�[v';3����_��*0Ǡ5qs�5{2鹙2�uׯ_=�|�T���4s`��X���{11�n��S�"����I7^1���8���i�N�BĀEy��Ivj�]���݋�LQR�Ɍb��Aqg�fn��<MV�rM��E\E��`~��(c趭����"�yC+39:^������7��X�1v��M�o��B�X���)� ��)����#(�o�
�G/�b��dq�#s���|����)x�*�?�7,%<>���(7~�"��> A�� ��{���QI}v`88�����j���S6^hþ���x��>�m-�M�k��ǥ���R����%������z�>k ��4�9�ƸZA�r&��[Sǂ3+��oՅ��J����nz9�ӚA_l�B����80D6�Xs$�h��FmS�K߆��":�J��'Yl��H�y�{����[�D������S�f���� v󋯰�/������O6������r�ʈ��1��b�
�XV�,P�]s�{���I�n�0��SK