XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����|!�o�l�mwT�`�I�xV? �x����*�7�m_%c �+�$;��K��h�ѩ�����qܒ#"�$�|̜��~�E�0)����[�UjD2�G�X�;����g�^4s������T��m�8@�iu�V���eư)���=���K��Z3�c�8����q�X��s4zh����!���DR�ӵ��@%t<�Q�� R܋��M��
��f�����#��ҕ�w
X��*6��Ӱ1�d����Y��<a�#أݣ+N�rw�_� ��Tz!l�������,�Қr\�4KIQ]8ɌK���8sٷ9@��Ev�3�9��ǖG=�j����2`�k��*��;/�}o�?���HG.�	���w<g�"bWKˤu��s���X"�ya6k�!V�O#���{�O�56��I�i�S7�_�f�IC� 3N�����U"��2&�d��^L[2�%\�1&��7�,c4\�<�*S�̫#�δ�"S#���(Ѯ������B���� }8oF*ʛ�0߸4�����?�����V+K��SW`
�y��K�w�'p��d���~�z�l~�\	:�S�[�i5h�dh����]�8$`�w�&��8�r�s����E����l������J�W��JjOvݍd�{3X����"_#�.�c\
�2f�?\�}q�wp�O@�����9_��1�Gk'�8m&t枋�����6��Aۛ.�ܱ��=��Rz�`�ђ�N������6k�-lFMr�#�b'I'�XlxVHYEB    fa00    2520X�I�ǱDUظ�x�p��̵��flF5����{c���
��A���8g4�A��r�i�b��TҨ���֚k>֟�B��|��>���.�&��2�P�*�M�y}��ԝ�{ah��!�����	է��4�����/g
ol6)��Sf�G�N�
��  )(�0���ɘ^'�#o��4�n�$%6���2�G7K��g6O�m����}��_�r×uC*do[� ֓#�Ű̶� E���9����a�7d#]i��??�^�g����t�>��g�T[G��np�_�D���f
�ΕR�!��83�gJx%ѷ'<�{u����G����p��Z^���YHk6{Zt99�����v�w���zC��]}
�����d|;A��6��&�,�K���8}pT�FKk�Պq��^���c��.�b�o�Y�3&θ��9&�H�<m�Nl��/�c�k80��0���uA5�����>��X-*��,�Mܯ{�|��\���#�?�h{ DҤ�9\�]�E�����*�ϴ��s��\`[���,>L�Si)i,�a��A�r]���}����I�:�m.����S�}��\����$T�_���`��=l�3U9�Î��%~I��z9#��p���O��)�계tl�� �9��c�����8X�"He�@�=��Y�c{;�}��6jT�a{h}Yh$���oʋ�2%�0
�_N��Tb@H�ۡ��;�p�Ho�l�`v!"u�ݺ��G��h��pں�&�A��\~���>KU����39�z/Z|�!	ꜮS%ˣ�4PO�R4�uL`�?j��1uǺ�z�\������|×�{cw�Wݓ$���>����iu د&�������m���7<b^�r�{�Sd��}*^��.5|�,�L3�J*�;�B�kT���zW �����Z��5�V�L�$�?pe��尊j��U�]̋�@ 4]�Y�0�R��U pͷ_���;�!�S���e��~�����{�|0c�Z�q���?��(�s�5s,*��T��D(��߮f���Cf[ز2Z�B!�Q�E���}UGE��QտC]�X�kSQ�?�=�xb@Gk[���L�T*�+Xp�Sr~V6�T�PP3	#� �E�r����xVp�5�9#�Vė&��� �?��wg���������`����N��¶�Ym�����H�B����6n��fN{L�Vi��\E<���D˖ln���e��x%D�+�P^Q�7�͉�t�|~��-X˙�̎�]��;��\�����F�2̰"�-�'�����2
�fl�{s��ӂx�Yd�+w<4iv�����j�pm���W������Ɩ���+æ_��f��~�y��B�����߁�)T�^F"�,ܜ�5E���a�D��������4�$I���_=���+c<��X;	X~唼�WV|�� C���Ʌ'��NV&]��qh�N����c�/�("��I�De����rà�;�U��`hez�"Z&Dl���>���Qꮣ7��A���p�3�NY~5�_�<�/ǣ�P}R��Ż;/g���H���R�{KҬ<ĉ��_�Q�d6}BA� ��v�)W�on�sK=;B�J�oh94�v�gg�ڵ�=����!8s/n�)~o]FN���*[���(�U��Wj7M���KX<ؽ����?��A����B4�~fԮ�u��$t�K sC��v ��O��d9IɘH�-6手zl���S���Q�����dޖ?0K�6`�Y�W��_Y^+�ε��U��ӊ��y���Q%Y$�mA(~m{��[�M�h-�Uj|k5[��)�|H�i��{"�u�ܾ���X��ݣDX��˅11N����)򅅋��N03�.-.�z��N�:ad2�Q�?./��3vH�YÏt�fF� �<�l�8Ux+L��gFcu3��1�C�J&��$u�Ba|����(�^a`l�,w���H�鰶�={�x�r�~)���"A��ӳA��;F���5|���_SS�Eo;�.�=
�~,����P]���6�YÂ�]M�tM�U���qnj����W�������҈q�͠mx>v�LW[��x��{�g)@A�8������ʹmP`??��e���<�������Z�U�����'�������wc�zEۘ$�a�G
k��*���:���n�R#��OaC[�'��=Z�����N�X�k�ᝥ�ȍ���ǧİ@[p�)|C���٩Qb���9.�~y/����C��g���S<]��)����߭�F� ��^vNR�5��L���&s6���\J���]��?�ƕ����j��ȀJ�ⶹ��J���h�m������糵 벇5�̉���6���%��ucǶ��8r�ǽ�SN8���B6:�|���Y*��M=Rvy�?7'P�Ls��w�����mI��]�f�Ѧ���8�ez��0�M�]�6�����Lα��i���*d9��?,��L~c�2���aS$��� �bH`��h!F�!��C�X�oaPJZ�:�Og+ J�lϒ��P��B̓�0�4D��@�ϵ0F��
w��n�
�M����;K�/��M�*W%��T��!��EL'H�oTQ� �o&46;t/��n4���ef�`���us���~�BD���Yu���V2��.��&�jPO%�ə�N�N��);~p��6-���������@|��I�<���3���b�l1 �ý����e%ܡ��3<��M��A%q�gaE��Q�Y�$��ߙ��w`{v3�Xh�}��s����~Ɲ�
���m9q�sЅ1 �����o� ��V)����q�yE��l6�+���c�A��X�\�h��/"��X�X��#ʖC�ߐ�WӉt���[A�'��&���5�cI�kfV0R�g��*׃
�*H�{G�G� DO6�����G$R��"�$�|8��J˸�V�T#n��%.Ј��>`����1;|�ވ����L��g�eXP�?'� �J5O�_���Dg:��K��*&(�iћ����wh<�&�Ũ�˯ﵚx����R���^������Cֻߪ�m�U��w)8F��Z��+���Q�VB�z�&vK*���e������x�g� d2�y4gb?eR���m�N߬���F��c����v����^-~�	�)�i[����
�|�O�"���|�_�&���^��+���C8�vLѩ-�m��R�,ƍ�4��IQ����uM&<�D�_U�X	 oD�D�@�I H�(�=�0�r�ŌוH�3��͕��B�3X9_i;~�+j�aF���Z�(-l7�;u�hQ�:v����IE�S΅���9v1@�Z��ׄ�)����c<�ӽpߟ�@��y L8�,�>���ջ���r^��{���[�N
�q� v\
��y�TmK�
�B�Ч"uB�%���ΎL9fqc�������w+\ݾ_uj������^,���3���4`�Rт�(`4����n� ��i;}T�5��wW�,��0	j(��2���z�_(��
=S�M��{~Rm���gP�XA��f�F����$ȍ�t���s���I�^�!�;�.�U�/"�l 8�|��������P�,|���F�y=�j�A�s�sP.W����b�Zɒ6�{+@�E- t<S`
J���4J񌜷/�n:ޛ�0��q���'��{�~o���K�7����{�CvK��at@��������)j:d��u� ��1"��R��օ5oF�y�� ��$u����M��Ov`��?��*�+�Fⲵ6-{p�:)�{�S�u	N[�,����ܝ:���j��_�<Ў/��e�~���hG+̾7]2^���&a�/'Ⱥ�^S9(��r�py�p����f0��n���+$��R�׊+�r$T��Xσ��kj�u߆���q��%�z�\n���Ew.9R;�'ν������qA"�7�1�y�(hF��A�qE	��:�}�2Ϋ���_�ls�A������B�����grL����� �)z�	7�h
�R�=S̍q���O���:�Y'���B��B��)
K��[��M��u�n3vbzU@��R�fg�ᬁ̟�l�������h]��`���S8Ƌ��D�\^��m�%��݈�߱O�f���xyƄr���{����E~�HG�u�9�$'�q��xF���!H�X2�gx����Ր=P�Ӯ1U�nҒ�j�C�Z8�U�~|�hfȑ~-T��`�۝bP1��F�6���3)&��0�#��'aw�M'R�Vo�!�=*<DJ!����3�M+*9z��_��j�'���X2>����U5��<�xnV��r5���o���ݑb�\Ҍg,�\�&&ԞM�m}�
mSȬ�i���32�AJ�$��\^똞X�l��f���NͪR��U/9��ў���-.7Ei���0�
�x���Z�=��F�H�5��jڄ��(R���yܖCy���Ѱ��`����Bv���UV����59��]>��y�K����Ҡb�?�T\��X�[2
@�:������Z�m#5U��%��-�ʦ�#�C1��N��G�5�ˠM(�r�|?�q��&\̀݅P���dmz�h�C�`���=�1��T���j���v�-B��6�EIs6���֛k�rw�닽:����f>����'�gl#�����  D�#�*V�V�;����݉�V
��=^`uH�߆�/7��� '���Yw��žX/ɛ���L�X:1�)X?�|�
���o����ڽ�����P�*삛�;���snX=W��Ufś��C�*�)����.b{���I�҈��kR�S&
/(l�l�}=V�v��M�n���ԏb��1W,93�=��zL==.�p�g��p�}E�4��X�e��T��'���ڍ<�C#y4��A�-���|��hͫ�rLD=)��9�_���v�w�U�/}�V�|�y|ơɞ�+*����6ج	����z�z~�r}(���ن=���B�d;�lk�)�.V���a]�����E��?��z9xT$9,ɳl�Ӌw�4�K�� Ve#H&���*3ыngI��>&�O,E��K���L��$cW���<ᛮk\M;�wѪ�m� �����}�p0^�GE}�9Wc���	�c6_c��u�r)�B����������#:a�!fGV�X��u�Q�*�y�BS��QU��vHw�)_��mu��Ez�X��Ŷ��5���v��*�`]��
�E�S]@��"��7����~l [Ï�/�N����6;$��V~�#T R�9J��y�Z���J�%'�UK�"{)�U����+ؑ�r(CBH�G�ȩ����<��i���iЀS�'�aaH�ld��Xc�z!�F۳l���Κ
!y����4b`b��Eƅ)q4�G��h��"<n$�4�Ñ<A���íݲh�&:�������a�1ȥ�/�熓k����3cq������o{ր֜�k��趷͔��F�*sP��b8���LP��4rt_1͊/r��c��f��@���9mCl!Z<я�6���Ǜ��9�UL&�(��[����V�M��ww�G���l��]#�Δ��"&��r����Pn�b�b@�/�HAu[��y��}�mm�a�7uR��ě~0o��s՗���V�|�pI�H��?T�y�~��k&��*�m��r����sF�W͑_6|��#gK�l�0R�O�e�v-"�G�s���ED�Oa세�{r�jLԈ�,�>�Զ�m+9Z`�����/���֧�F��e�?�4m^�H��7u���H�-HL�"�4~��-�PD�:b����&���Gl�M�2VLG�����h�݉j���H�]�R�S�>.cTUٕ�`�JAv�3yrm���}tz٦��S�Կ��j&��Y��x��m�����֠��q��m�:4g��I���@�O���e�Q���8�̉eUu`�Q��e��>:�����Ej���v1@�)_�Lǐ���������$�z���ѵ��|��m��w�,�O�\*�#(u��&Z�9]�(�Z퇷zu�� K�>��h��g����C�pb�Y�nl0��(D0��#��J���,�3�FNO#"���qq'��IO$7m���xC��@*�����gj=� �O�1�Êp�$��KDÌ�`0^�G8����Aj�B�.\,,]�缃����i�W)��e!s��2�|�(E�@	k%|��G��.1�WP��dBS)"%�:��Dc��Q��*�
� X����+�BD�C𴋢9������֣x+s���e�;[{|F��dc�=@�`��qx��zU�|ƽ�4��f�edHF���D=��7�]oZ(8V��n2 �P�b��MR��r>$Mj�������p'�h�R����kRe(%Sj�Rc��)�q����b����Dqt��V�J��[�i�� W�LQ�lM����3��W3���YL'v� i3d-A�}�i*�������h/�> ,b����-;���M��m���Dd{Ǒ�[���ܰ� �}s�4�y#�:w/,�@�ȓ�1Xb�;oo�;��}S����\�Ŵhxn���O��<�2E�dj�U�x��j��6�B�F�k��f0�9��r�7���lgo���]$J�M}�*� 8�Z22ԧ�+���-���)Vem~Ƕ��P}7��h�J�v6nƢV��x��z���ʗ)�ddp��L����ණ�1�Gk���Z�]/�E��mR�V�6*_]nz�]�႟C<��ݼ� ߁aeb���*;cq�����8��Kgw�!�0b��lb���.$�v�z��F�bA\����X�t@[��CL�U
����D�+��f��ӱfڸ�'���I��y?i@8_O���l`��p���-~,�ɇ�����TQ��H���M����(C_�V�tf��ځ��$)�Jަ� bB(��1��D�hj���S��9�ƗW�`%T���"n����[τ+��/n�]��Y�5���6���nmݙ#�r'��M`� �Rv~ɯ����=<N/�I��W����ҹ���N�9I؎+�$.J4p�����B�ż����I��"�|qklO�3���(C'2����]��hU).����T�w����i�K|��HZ��"����GsNR(�
��YHւ�H G�4/V�(\�5����;d�J���,UR�r��.�_\u��C4~y�\�߬A`� �,L2D_�y	�^J����lr~��^@|	���=<���iҧa�Z��Q��.}������V��C#�?�'���~H���Q��Kd����du%������ۓ�O��(7�3:��N؉�w�C��	�E�+�̚t�s��Ls��[��N���%��Z�3�{�	߹9NU��?My�!���O	9+:0�������R���zge�J�h�l�֊�1*頬G?�m<�O�S��s�`�Y18��H��Ea����<g�~!�r}v0��Y3٤����ן�b�����A���/&I���k�Ù�e�n��lC:��f��~s=6<ؔ���@�Ss�v7ל��ʑ��$�LO�뼷c͉�5p)��(��������0�� QQea\Ҵ.Dn�2�H:R0�W�Gd��g��-���Ɛ[�Q����ˊ8��cG h��p�1��y�mᬖ}���D0sc2����nV����{����]S]��S��\i(qux���I���`�J�s�f�
G=�`�{���S�����$�zj̘!���7t�B�y|T�k\B��	(q�	"M��7	*G���&X�~��E_�ּ�Yg���8�j��t��h�� (�G+�v��U	�>�I�����37��w�"0t�bN�n��C����o��/$;�͵�F��U,r
=g�����:� TК Bڄ"9����1���@!spvd_�EF�%"јXS 5[�5��c�قgo�!����=�=�R4�$�4}� �T�r(.{^ ��E��+�MkD�Q.	��ho0�d�>N[��@�	�ӯ��r{q�~�6��M��"@�)�GIiB�DT*�#U�
YO�|�˶U�G<���v7)���o]���J�W����>��yR˯v�	��p��k��VP�@���M�[)M�����TN��~8P��Q&�Z�>�Ѽ*z��u��;<D�Q������u�����CFjH������4h-"�?>��K�@)>��UN ��?˼�f8��KW%�u!�{ԇ�-��#m��O�j=�=ܠm�*!� �Mɘ��~���!��C��t�NQKH�n�l��U�.i��6e��%~��F_¿�����{��D�'��V���Ҳ�Dv�
�_��������v��Y2!���ьY��Y�5�,���"U��	H��~�ٹ4��i��|����n��M�'�wqv���t�Q�(y���s����Z�.Bd�N�?�F��-�jK�_q�J�8R�V�2vg�p���,O�Y��� V47���X�l_�^6̥���
R�����������k�[�Y��si��Р��K��1c<�iS�s�?I��g;V�����k>M�����e�7��c�p�x��*l_�7��RL�L��:dB"6�z�o�15�����ড]܊]����a����)$n��U�ŏc4����]y���*�$1y<b�m�'�-��ސ��6��*sf�r��jSBj�B����5p���M�(d�Ge�$��l�1���B pW�Ƈml�au�O�W�J��R�K+&��9�n��0�f�)�T`����8�0�8'�4��.�?s��e�����U�
B�`�ža`���y)��@sR������f�<�ͣ;Y!��d�p�`n�ы���z����o��o:j1j�L��"��a����ɏ NE��L:�ӤP6!}¤��lAb�-@��On��@.���Ŧ1fj���NƗL8n����4�9��?1�QA��-S�*�4<���I��.J��H�O��Pz�h3�o?�{#A�za-���ǘ΀ig����U���:LsGo�)�J�������[�mZ�Q`�1����yü���`Aj�0G��ݺ*>��`�������ޅ��|N���fע<�/=��������"S�r�D��α�sD �)���*�Q��F���d���g�8��f�'�,~���C�^�N�P	�DӋr� d�Ţ��	��}�e2�?Qμ`l=�@H2�e�h/ŐRp���o1���OT[3�K16���F55��JNw��9���L�w���g�BY�*Ai�_��d�52�#L���+���W���:�-qZOb�0XlxVHYEB    fa00    13e0�p�ʒo0~�c	]�sb �(���R礴�O��ē�Ҙ�9�z� O@��z?XKC����Vg�*N��M�v䗇��Qp�V��aC�2
'gav\�����Vϛ�=�?�5#��G=���8�Z�R+��#h��g�����B.J�Q��y��5A�����аHش_�;��Q��VL�v���[L4F�?�տτ4�+���W��W��/��'��A�ʵSo����K� ��� �E��p��NTK��UE�9�/�q���[m���ݰ߇�e|b�Ξ�K_���o�^	a�{��n\�6����IA�I$]�©g���Kn�2n�hW�߀ƖX&�Kű��B�!�_6F� �,;&m��IÉ�m�N6A��U��kkB��}\��A��h!h�YA�J��"���߸2��Z��0L�GZ�DW�e��E_س�vI����fY�&RϗSJ��6�9=ʹ] +U�'J��{п�ഞ�#뢢DX<8�@���D0�3���I�p����꣘�VŻ�U{�[�T�D�>EF㻋�K��i̞SDم�W���K/:"�&��#�����I�����n� >?9��64#FS�U�w�]:k&�D?5Ml�h-2���P�,ǣ�J���ܟ�e�R��3~P	�������7�}��X�0>�������W&�f`q`��4d�Ħ	���oPߍ��pT!G�C�$��[��pt��8+7 
��	*pA�Ѻ#��Ձk֭^G�ށ�3��W�__\w_A�Ʋ�r;L���ȂIBŌ��J�Ϡ�1 �ẖU����c�Po?��Q?��o�����s�f����u�z��`}p+hss�_:��ۙ(?���fYP���H�=�%.�{�X��)�}��jK�g�.�	�{�#Mۤdʛ��ws�çY ��_hqJ�hə����ΞK�L\-j(�Z�x}��6�H��>�%B�~Nʑ��}��4M�ֱ�7�7Y��r�s���ι� Ӷ�&��N�
�b���W?�X}x�hL��ߚ佥G��>4��e��Y
�G8�)����}�>�����.���5k"�)J��Y�N�!<����鯀;#�~��Wn�	ٷ�D��ʐ5�������9e��t��k��:��o�D�$r�p|����}�C���-�[�I?p��	��ƨTa���;�.Dɷ�C4���qu@��t5�0c�KZ���0�a�o'x	��U:��^�g�UHxLOp��2�}�����;8�dq�k���,+�����2ؕ���u�1��Ls���7ST�e�oہG��W���R���}��mP�����]��^��{'C��%��L��o� �п-_2ܯ�Y�� �ZU�]A<����f�+�s]>e��v���;gqJ�%�jfzc)�#.�j�8z�P|%g�������.\��$�1j���it��ө�$�f��2��t8U	-��L)���*5 �;Q���'�5�)	��R�;jMY�<X�ɾ(_�d�	�r1��\���sB��ڹC���~�x)�R�j*+��oU3�j�c=*D��ێ�ZBM�v�X���W����ٓ��H'�a�.&�$	ې�e�?�qfh��v��uJ ��;X�p�~x�\o>�!�����oF۬aVO>�D~=/��D�+��D�f�d<��b�>ߎ�Q�����������s�e�;���p�ŭ{�y�߈�1/'nRG�F���Qr����Ɠ�7��J&zj���2��� ��
�*���:wB�+�]o��p�rH��0lG01��c���?�����|��z�J�����H'Qx��B�� ��z>/�9���e���	T�:u�Ce���>n�fh�	�|JQ8�Ra���P�}͠�^yk�*Ke�vn���L�+�ɡ�m��[��O�!d��s�$e-���' ���HLO��!�8��Rg�N�@��E!�?A��U�OW� �J��#��� �5�´ȴ��c������.�@8H^���Gc���I��R1|FԩPd�.��xA���Ez6VG2���*F�_�(��b:w)�I	����~b���Ul��WE�������p�W��ר��v���������*?I�uL[��s�X�{�&~����-���Q��tx���)��qM-6%�@�m�]��2�N"��ki�@�[^�1減nTԄ��x�:����f++{,�ύ=֯�>_�����=�#
_�q�������C�ο�­[}����د�/������Ϥ�C��rYS���Hӛ�ÿ�ע[	���UI_�I/7��x��Ҙ�'�JHļy[!�}���w3���
|���w0��4K����+��!gqG1^�:C��-�X/��nߤAQJu�|����k�.���G>A�MnK;ug����ϰ�[1���8���ۋ��^!m����;�����<���ǡ`��D�1�}�p�Z�˕�9��Ɣ��:"B��`��ǘ���_v��a\D9ZUu{S�8�%�>Hq�;<<�<)����ҕn�;��铲〕~]�á�>��Ϲ�}`;Ͽ�蝦�1��4=�(8~%	�y���ŋ�.��]2s�;O}�oL�u^j/�ώe
��Km�ʷ�U���Զ!�8-B��Z �o^,�
���}��7"���@��q�2�p��E��E�@���u�q>U��ʀ,�Ѝ�������x�'m)���7M�4�s����||�س�|; �d����s�������"� q���i�=ۨ�*�ۏ;-�������$}Qsu��t��V���uyC8+X������(���}����t椆���V��� nT#���ρI�/@;��H��3�ǚ�@v����X>Z��D�\���ґU����bI�)��7���F4+Е��:�L3�g����\/ŕ1�'77�'͌xΑ&����x�t_ ���k7��tbg������XX���4So�]]4�1��%�Ri�ف�*�	ybRq�U8Z�v��#i�����v�2rL?�#�xϊ�6*GF]g�gƑ_�kkN�����=I��*>���i �5�����T/����9����PQw���]�;�
�%�vMג���ev�t�ݔ���e��8Y��(��S5��f/_��1��+z�Z�`��S�S�=2�L�)/4�J�;�Z��aU�G�{�AŁ�3��Nq����H�Al��H�{H���ba�����H�~k	o�l La����ǵ��,��Ec[d���I�
��
�x�hOȅ�5F��S���T<�}�1m�Z�&�=�o����9Y��Q�&D篕���dH^ҟ&J5���_���
%k�j�A�SE�M�5=S��S�/B�
>�8�D�NC����'`�ㆴ�U<���p[���f���!� !�.�YH���n��*�=т�@�5D�U3���V?�M5>J�歧��x�w`^�(Z�LG3�+͉��Y����2����Zs����;��I��^�#���d���+'jЅ�{T��.��eo�9��;m���3����H�����W�ŭ�E:�j�%��L��X��@�p���o��r��Y��EȊ���d��!S3��]�F��	�׃l�A�byE�����߇��M���帾��,�OϮnn�[� ��!���*�@���qd%q<�"#���3e3=��B�Dc��H��9{S�����|sD�V�;��&�s�no@GW�1�3/e�Uӱ)��b���x7�Z.�M� >N`o�'zM)�!�ݻ>Ͽ;0�h�I����uU�)�"�v��A�� 8�	���AO36��}z =c�f�ݲ,�z�ܰ�C�􍎝�D��0�r0Py��N�/�;Ϝ��A�c���'�݊"-���h�쏓'�"����A��uL�k�Y�?����[2�'�񟂥}�0�"J9B��s}
ڏ2r���̄�~�e�B���T�0̍�i.V��10��9����S}el�����\m����7B���)��j��l���zS���ڷg'S�v�5o��F-��>_�ǏO��M���E^��	hg�Xb�a��EܴWq2)F��؋�bԈ7U�a���>2���N���i:�NqP�aFg^��p�Z�b'ӥ�d���e�{��c��b[8G�=.&��A�ll��U�q���\i�蛬v�ճ�����w�m�_��l�VamD��T��֎�@O���	.�����s�"�[�r�*du�=�����/!�"['�ɥC ����R�~��C���o�4�=-ߑ
�8�?�Kg̛3�^O����u�2f��2�83��S���Ӡz��?z�֛p]���
n	���dj��OU�����?���8Ց����9�LGZW���:������J��X�Qs�Ng���-!���d�S�<J�B���*��(P��36�J��|�ZP-�1�a�^"���zձ�a�r�O���02��j�6��LÍ��ń
�t���	�nѧ]��%�ƆJ���4'��2�pr�r6���5�OY~I�k{oc(s#.�?�
�{�BȾ���W�0S��z��b��_*t��.h��0箛1@�#���6�Vֺ��F��l1[�}��c�T��v�!E�SW�Ӆ7��7Zݙ*�&�t��@h��O�����t$�%�%��,��T��m���:�r��֤������Q���W䦗i	�P���e�\���l)�6C�S&kfqH���/Y`(}�)i�HU^A���5Xs=4z�ZΕ��H�:�J?4,�^ ��d�M�e���#����R��)�h
��7H�j/���60�Ãc4Jc\��i+ońQڠ���Xqy���zD��!!���h����d���k����`����pτI��[Ϝ����ăBAH2V���A���z@���y�;�U������Z��}b5.5��:�	6Q��$T�>QZ+�@ڠ�n�Ƒ��l#A=q�po�X/���ܑ����XlxVHYEB    fa00    17803�%���30�����_��U4@�(���;�:�P���#���%������P���6a�w�
j��/�������s]���pi����̬S}�h�ѬU��/3�Ձ��:�ޅ��*� �K?����!,�b.�#��F���-���,��5%w���Ԋ}(����o�/������7���CfA�Y���D�d��:���D��V�]j�V;���Q�:���秓���s2�#ý�2�lvr��`Þ>��v`!s��,]��w(+?@�������"FU�׻�7#.u�{9�8h�i�p)&Э5���\�7�?�cSɘ$����dBm���D��'6�`��n$���	��V��7���:s��nk�BLʣ��`̷aN�͝��N�y�ѷ�a�)H/x�{�����A�Y�D��������K���F�:L����G�KP�>!�~���F�]�K�id�>{�!��.0�Rwp��n�Z&-�/1������(�8H��/3)��).w��s�Ex&$p6ծ����n�o��i�}�X�
�2:ʟ�o?�w5i�m�l��ϛ�0"BT��УK�[(�vy�Á�Zĵu������puhm�g���~��Y�d\�����'U撦������`���,�E�%���� ~�8����Ղj��]��N���Fޭ������bS<3Y9//�����I�5���_B�Wiտ}Q2��8�_��<��:����<������ޤ�3���C��/�x��vZ����.�w�b�D�ÓC�g�D�G׸���W�*�����mP)Ή��	([����7"�{�lE�GK�R��'�B�	�H��V��'\����=�I6��m��>K)�#�OlE�n)n��� 4�B���}�����T=�}a��35���P`�	���Δ���Y���-��ꕜP��6w�m��6�W'��{j����5
2"ߚ� �6���$��� ����}�/�ڦ�]��#k��K!q�}#���s��JЈP@E�n|�4S��m�K��􁄃V�z��v5�H�X�{Sp�����[�!�Y�3����b�y�U.��E���툚X�&�ҏ5�;p��H:�{i$�V�i�Ak�Y����|�b����%^u\��Ӧ������⑳5�e���8x�����d��P9+��(b�����jeh�h�����@y�O/�BK�<���.�DUW��4�@`����m8W��mN��h��<��';K��уۈ��Y�G"��S[N�*�S\z�Ѫ�s˿Z����#U��� qj�3�Rw�+�[���u����Է�<��8:�|�
�u�H`��N��*�ں��n�#-��6��ēZ�K@<���u�H�݆GI#y}���^gM���¾
��7[�l�q'tIU�yȍ��7L�a���t=��(���T�p%�I�^�����)K�T2յ?]'V��
p?D�`�C�(N��B������ӷ�<��8�ZR�F�+��' �	�� �I��_lP�x��s�����EUi���|x�*6R¦5iчUqkf����RUAo:b�K�F���1x��*9���Б�2
�a7y�ķ��C���H����b6�!��6���ɜ�������c��7��O�=�������O��X�*i����7?\�*�U��u���#&~���#>��i��-#���K����	6;(trL���N)*�aT�΋�������P��"幣O��.��s���7O���x�j�	?���zn����'�j	�`��2���O�u�>��ɧ����[�F|�rw�0��u��s�H����d���Ymfg1�067�0�tB�<��X]�7::�BJx�_���[��MO����ܲ� �|�e�>�+c6�*�5�� �� <�}�D���E�s~	�����妖(?ظ�@C�T��~�JqL���-i����2��q�X�
�3�.�>bҜZ:f^�'�wVy'�S-^�z"�i~��ve�̀�����H�.�}�"S���M4�L\gC��u�3а�	���A�R���G``Uzs��'�;�K�?�Nx�?�T{�_�f2$�_<�su�[X���B�L������T��,���ї�Mjp8���]S��Uo���-��#)�ɸ������xo�ځn�W����4oOؖ]&��������ŷ]S�n?vW�&ɬ6��[u�X��8�~S՞uF�
��d{��e��	ݥZ�0����j�~�f��BnuwXp �j�2pfJ�$�bz�!��Ǒ���n,܆MI�M���#I���j�9��%I��k�#:���<�Qd�q����,����vB�j��U5����Y,&�d�x0�4yd�=%#hU�!����v�+��A��{��bV�~]a��e���jV�dgFQ�xk�n��:q����i8U۔�c�X�e_�Zx��7 ���A����"�r����4�>����*D$��I��1����弭q]�i��%�;��ki:ny��^7;;B���n��r�-S��6Y]�|&�#�C�wc�d�%?.ļ�5y3�Z�kL�g�#��$i�r��K���L%s'"�����e�a>�M�E{2p�1]�ne�@���VE�6J��i4,ۢ�e@�;�L�X�^d'�~7�ۼ>�O���8�~g�P��w��
��QC�G�ǔ�����[D�`B��c6��M�zN֤ӓ- D�p~�=������1[�%*Mb�tJ��7u��;�-ݵo1��oʿ�"��T@D%�l=�e��B�B�U����]M���OA%X�G�ݎ�%�u~�!p�l�*vS��uNFY�����d����aPk�	�|�L�~��;�[c�Gڋ�K�F� ;?�=M=s�<МmY��N.I,e��Ks����ο�1��k�<_��+��	)��9�S(����?�D�\��c�:;�U�V\��v$���t�-����D#}�B9�=��]<�_�Ve7�;�Q�_Tǉ���G�Y��pIl�D����0��b%��{[&%PFȫ<�c�3cV��Y�@���.s���#к
;�9�$z��
�JL9�_Vh�/�ig�#��b�e���{ť�x*�d�co"Q�53^�|�:�(��Y�*�І�eM[*��G�}H��>J32zin4!��B~`Gx��j!U�B�>�{�NX�W�-���:��?�MDe��8]��A$����e(]�� &m�*+��PO��ج�j:�Rȁt�<�v�S���8!opb�����M�X�q��FR�6�Y������}����Ka&�,;���I�n�܇"�>�z���w�Ǧ�3Ȉ���ÑC��#^uG��0U
��g1P��$qg��=�y΃�9�y|�"*��hD��fL�S+�)ö�E +�-�xwbH\Cv��Dq��բ��^DAq��
�>aؾ��'�=,7�Z���FE���j�a�$>�*�*T� ��[��{X�<�`R����Z��N◙b��H�R�:�5�T�By����u<W���_<�B��g�C�$z4�§Y�בּ�å����4�Oָۚ��¤�o�� �Z��}Â��g��'#�o����'�W��d1[�B ��Z�g�ն��FyG8i�H��4�5F���]����"�����BKvn_v�}܀>*a����5"C�S�m����\�1��?�:��O���_%Xׂ�r���f�ק&�WΨ�K��es��� ��ר��L�"J��6S�F@���� +���@2����8.`8�|'i��ߴ���ј�0Y�Y�dAULc�@��=ut��B�j��1��6^�+�ӖzYz-ψ^��]\k�&{T�0X�N��0��ȩ�R_d"G]r՗�v���9��K<k(w���"z�u�.�+�Ւ���B�t��/���*��,SB�3lʯ�}�Zs��.���{ߥ( $�R"6�a��/ē}O�Í �Z&5O�}\C�X��B"!�LP���~ܹb���0��CC(�!@��F�w��N@-�����a���$�2-N�J��R��� ��v]�!4��2Q[�dx���k`k��AB�<kXap,�T��.��|�8�r�=�<���g�Σ4��REoHfc��.ǌ=3 �z�,z�H�y�\1�����ka��x�#�U�� ���\��X�>y��OqXf��y��-�A��,�L�pd��h���5���
���taj��h"ʼj�l�N�ϳy��͊����P2r�-$Ŀ����@�w�Tl}1��D���s��̒0��A�
p�^���D����~�(�����p��{���E�NVQy�<˕��H�р���ۇ(��8��>�" ΄B�ĺ�!���P��V'c���Ӭ�;��=��}"�M#�U�ѳP��'x��H����z�yRk4R.��6�;Ӌ7��.'g>rl=�� ��/����6�%FÄ�7J�����P�t����S�w����N������e���
 �̡#0�-햃��T�]��q)�p��b�X3�.��Иjbc�~�'��ʚ����V�l��!:M��,�x@91|=��PW�AVE������hC�.`�hvI��a<ФD*kp���2?�E<������由����.EM���_ ��7�̂�����	���#ecfA��C�d�ě�����!p��$pڤ��Si0�l��y�	_5�����n��5�A���V	`��w�
�©j<p�9>�@�.�r^�D��r�i�:K�������l~���_7ݲ�/��;س)8]���E�qةA�:�՝���y�=�����4�G�<�RX-��h^���q�W�S�n�Hg�<k��t���qn^��W�R���o�CX6�?�yO�<�Sad$��>�aN^cI�ILX{k� �Xe��n	Jt�-�K�(�gj��tJr��4��!�P�$I,^F�FPl�=џ6_=�W��O�!�D覉��nC�v�P�0����k��#�ۚ��?ǚ��ߥ��*��9U��*+���z�ڮ#}Z1�/m ��C�8�Oj2V�!^r'��C�!s�\{bU�/��ܣ9�3���_�c����t%��#�5�L�"�� L�v�.o�-y�$&1�*Z�Ix�Ao���y��G���Ρ��nk=kt�BRJ~s�f'�^�L���3Z����}����ؗ��%����+
���}x䏩����J{H���6wu�����5�X��IEf�(��@����������V�Ґ��zI��v<����V�ERz�3ҷ/-��� ,��c4����][�wVw
�;��%��x�G�z��=��/���l�R�%,�����Հ{^��-V�2Bw�;�8��p�jV��Q��I�?����M�;1X��y4�A���3��[o�����F�6dF|��MTU!>U^�֨�:"�M̩�=���v���lo+��o��&noL ��qD�d�E$]!�e��/h{;�m��S�]R�a�5�+}�7-�Gav���� ܨ&�c��wtf�ĭyƉ�ݕ��X)k��m�H(�2�!����77�$��4o==-lNb�d���f9 ��JUu�	͉�E?�~��n�(�PӀ��f�s�
�ߙ�A3��
w����
�������[��cTܹ%��%
k>�w?H��p=t6j�nh�jr0��Q�a-�9��F{�I#���㇢V�l[N��*<zh7��j���j~:Ns ���{{Krw�CO�,���5n`�4.f��"6]n>��#|} �	abiw>�x����NxC�ܛ�r��5��o���Q�m�
 ��ξ\�h��a���s�B/`H�/{��G( ;��c�^�O��}׵�;�/�D���d|[7���"x��[�Ly��Ϊ�*h�7J��-/F����/�Wm9�~[�3p��.1��l�m��Ǳ˭�XlxVHYEB    fa00    18a0}�4�C	f��z��)ώI&$��R�����d����^P�Ur;�=���4���n�9Ģ�۽%����_���&��A1�IU����_i����:��`�.��K���W�����i|��N(�R� �id�+�*�E��0�o@�*�r?�ECpG��hQ������3`8x�p��yd~j>�q���e-")�řز�T_��y�O�o�_&v����&L]�Ք6�,
���C9N��g�ËZ�x�yo�� ҍS
��W�{�;�7�\uA`U;�/@��D_��A ��̾�n�����ٱ�%��W����?�3�Y��>�"t���-x�d��/����\_��@d<H��1��N��/|��gzS�ʲ�b�����Є5����3�x�2���h��Kgnm�^����b�;���|'6��pA�'�bH>�Vҳ%���3�]�S��eT�îOm�����4A�x�m(��8$����ptG'��c����G��
V1��
�d`$��!k���������6�"I�nz��bw�f���R��������W��<:(�h�&�1Ys�1n_�*�۬�*�_��s�N�!��a���oG`���bbi�ͫ)��C�8/Lhh�P�eH���ù����"�.k���1�^3Vu�p�%�A�˅����H���������In5����[*r#]X�ρ�VΔ"��A�%jI�����]���b<��W�+��E�!�L?ut�x"rY;˔
��nb����{:�����ME{]]}~�|c���N���D�E�%���X�e��p�`�[9���z�����&Oǩ�ބ�8�5X�2�����	f��ݗ��� ��{�*H�Jo�i;�s5���̾�g�6���X��1����/����r�3:I:� _�:�rTGH��� �q�A��r��#Ze�N�6D�g��O��E0���B���>cX�ls]̏]�|�is^Et����柸�0�����`	���\"�ze؏��HP���o9��xX����
 ��Z��pg��h �5�P���6D"+��۱����Y���t�L>c,!�߅o�Y/\%-�P���fuo�S��ST�c"L� �pBo���ǂVD�ۃ���<u�j�"���*��ds�`s�u ��w\���8-�W+����fu4�-Ż���44w6��(~�`�'稃u1}8�O��7D��k۷T~fa���}O���G�B��	$�*X��[d<��v�fK��.�8�UVG`t��ƃ̒I��(�N�7���&E��=����r�;���	���+ܝ�o���}��$t�!`Ϗtk2x��c�MT�?φ��*P߰��m�����9�\�2}	h4jErKF�x����*�|����]�&��Q_Zʪ�z>3�1�l�Fй��)ۛI�%�E��
И���*�2n�=ߥɒ�Ҷ\�i���Cz/������@�eS�(B1 ?��}9�y�-�G�Ӿ@7��l�-�7$��X` �������I���Գ�@�)���1�*�uJ� ����lX�|ۉ�R	�q���J�|a�m�u-�JM}�]䳔���ܤ�!����H��N�d��/XF��`H�ƀ�m��,��I��X��A�r3��vO���t��o���G���;Z�r+�B�R�Y�,�p:cd�BW����
m�bDȖ&�;2�&�q��@�,���`��c0h��כ0S�:�n���S���d��/�l5`'x�W�A?��]KI枣=N�Cu.���W�p�V�7���]Λ9h~v�v�<+ծ�6O� D?ۙ�W��������sb� 4�ف@b��=���I��,>k��c�b�����ܜ��XJ�B��_�Z�H���r�C��Fn�5T���[�\ �f�pȳ�W%��G_V�W�H����[�'�~ ��:�w<S���,�(�����A�T��Z�ľp*%�	�+�~"��:U��]���'򋵊.���b��`��P���H�W��9s���q�"7#LJ�MPZ �b|�	s\􃋝S�!�]��P��9q6EF|���.��ӗ?����O_?ՅH�4PE����Z�ZT���ꡗQ%�'�ZP)J�B7@�`)_>��и1�Я�@�P,�nk�j�l&T9u�7��j�	Nze�3{B��/�s�@�W �{B3[���qy�T�X�O&�f@,��w�M����\���-�b�����&~�&��i��h�� ��k�o;X<���V#� ;U�-ib.�T������L/�R���E�]`\���@�#IP�\i�k�vL��f'���F����R�&�o�9B�U򛳊ޮZ`�����'5]@����q����֝����Ё�0��}�k����a$���T���6�*�Rw ԎE�Ft5��>�ZWC|]�]��y����a{�*�������"K*�<Re��
5h��?�[;��ľm�8�d�:��?D�|E�h��jC'�x[�t@��}��{�dZ�חcX@�+���hg��#�-��<����e�|�"�v�f�����T�^��Z����mv$����4&�d���[ѷXN�VEsdt,��Z�@�N�ٳx+4�U�mc��Vy��X������e�u@�?[Ϋ0�I5^X��5�%���]٢c�JP+n?ih���~�p)��/���мVf;��F��1[�g)wx�R�9���p�SC%H�9jlc���.❦dL�d9�j��z^eQ��j�t灴��ފ��kQ���/9�(�P���j�,�h������^1�ڼ�9��f9��S�A���3��'���N.`�AE��I�3B���Y"�������"]ܮX���6�K2�')��gN�Գf�

G }�җ��6��������:!�s�閒���L<�\0%��C��ˍ��#�G�#�kF��U��nv%c���q6,�>���~�XA��O�:��i�5	���N͎��ʍct�zd���S9EJ��A�Y꽅T}�Q���6N',�����m�^y!m��|t-�qS�W0�� �ݵK�M�������w����O��f1��K�~{�s�m��9=�/�~��a����Ews8��
�ۉ��Y8��%K-�(�]�����r����)Ϲ��dB�W�~��)�Hş��W{l,g���j��x�䋛�0�R�Ft2۫`�Y����f���9c��uyk�'����4�Jt�5���yW�����n��g��rˎ̱�!=4B3Q(�/�1��Jc�����_ ��*��E"Z7�ͮ^��N�lŜ����M�2I�x�,a�fD��1Q-n�@Z�'>�h =���kܥk�WYjb���c�VD1�\��*����~ٲ��^��kRz�Z���@+!Y�ҩ����M�
���ø�,��Rq[�3�%	��rO��?��]}����~����h| ��n��G�&6��x�7�[�Z�St	 ��O�#t�zM��d}�3�� aZ�=M������oK���l��K�(��%)�U��R�Q��)��p�iW��1�,2�O�L�f1�|ݺ#�6��Ĭ5�&��-h��ב�d�_��rRn�p���t`���W����G�D�'T)%�ǹ?H�I[4���k�'�h��	��"M����gg���L��s�ĺ�/h���c�|� �)DYC��DqJ�Lq@U&�ge��N3�=�H�p�"lYk&�i�P�k�bY_ާK��8�����'��ƽy�
C�����zQG��U�������cڞ\���`~E)k�ӢqY���}I���ɨ������m���$�w�x7�N��#[`�g����=�9��.q *��Eb b��GK�����.��Oq���Ml$�@�!�q')�[&%��Vhn
^��|�%�0�N���9��tG�̠[�{y���*�����Ok��e�',;�(�����4�)�Ȫu��F�?��AM��������'0��;����rf3
et����w��v��ب���`W��I�Wԫ�p!���X� ��-�]��k�t8��#�O5U��g�߲��Eip�f��O��]���1GoaA���d�I���	fV}�7)bK�2�?
\`��ŀ �w�u�"%#�&B��,.������d�e�gf�V��T��I�ă�X$U���5��q�+I���A��Q?f�����N��8Ra��B魛n����d4��R�܋xG�����eo��D8u暙����D�����5���˙�9C=�8����NO"q��	2�\PO_,��!i��u1�� ���Gq|^�Y�{}����ye������2!`�`2������%�yԅ'r�̿��Ow��쬓s�f�����"*�T�6z8�ڬ���ʅg��ܛ����C��&�o���]������Կ��y`��|����}�!]]�L<K~�^^ ~��7�����(�����j�f��q�����Ţ���
Z��K��-�	��B �fĢ�vlR��h{�Z�!��ԫ���$� ����t��ȹ�x'$&���=���Ϥ7������(�ti�z�$���(+�Wd\���D_�-ʐ�_�<C��9�n��[��ڊ��;�'�]3!:trB��cNIf-�����3��L
��" ~`�7�dd�/ӠO���6Μ� ���)����E#�t���0F�� �^C~�9��*�(y�I�p@�?�}Us������Ҙ�S������6M�[^a1m�����P�a�vx�]��������9BHK6<�M_���A���0���4b���`�9�;��1��
Q��j��B��G�)�������Ϡ��B��"qL�Fq�ͽ''}�鳊���g�$U��^զm���Qt!�r� �x�>��}�����y7��mA�J��3�cՑf�
}��q#�V�0?
X\D��z�|��+ou�*��rvs��)����A�����eJ|$�To;��X@޷�)��?�gJ��a�I�����`Cz�c�����O���}�6��t�%�ߩA���X�(�a��қ2J��iu���\��@хw�z]R����*�E:[��2Z�ɠo��[��,�����^ڌB�^Po;��t�_�ؗڄ��M�X��x��>�"� ���ﷵ��QN^�:퉀�U��#��IlCﺤ������~ؽ�Ƅ�g��[����+�L�ER�fE(�)x�9���%���@�x���k�����]Q:>�-yB�qC��XJ���u�t�q�J�$�.���p��+��}E����4��&:��m�Pt��w��d#�r�P6����c�I+{p��0ƶ����f �	���5�wpT��F�������x�~�������|m�l�8��G{-Ge	'����_��H�_�{��68x�UO���nK[-��e��e������ì�猪QB(��""x>�~��h���Y�֔	f��*�{��{R �����m��J
��36�TW�N�	AqP�Q��]}��������޽�:f�$��y�M�|#�\T��<9���9B��'Z�uKO����#� ��Z{��M">���(�������?܍�ùE���.����o�BDeՁ��b!�=nb������H��Op��0���¦�Wۏ���yԛa]D�� �GC%��I�}&eu�a<Ly��-K��Ho�����o*	K��-�y��뭿o.�����V!m�[>i�:t)F��{VO�.�
s��Y��9?�湒G�� ZMQ_�M.�E@�C����c،��d��H��R=7�{~�w�2�k��A���_�"��8�����~6
>�Cf�T�Q$�pd[Q�M���/'"��f�����^M4�����q'��$�C�2�l�3��0m�'2[�@�M��0�)l�GK��K����/�-�~*9�Myj�Y,v&w2B����I�'��Z[�����t�=�{�-py���*�:��Ra�˃/��f���(nW��]��M�f,�J�?����M�UX��O���қ����{Xq��q8�����"C>�3����;�������	\[[�_�w�*�/�r)/0��ԙ>�/3#"M� \TX�������1:~�Ԁ]�mHK��|>�Q��V�,5��ᩭ.��2��,���!9��-��'~H�z����_۽Ԓ]g�|/��S�/z���^���|�@���4"�p&�t��L�?˪-Jک��dbXlxVHYEB    fa00    1200���"��"w���U��#���g�W;5�`G)�f���O����ڗ*zϐB[��ߤ��I����)ާ�O�+� w\�C�}�et�$��&	Vݺ:Y���2{��Ss( �c���5�O��)+|�\�bD	K�;@����sKJ*3���S*�@�2������x g.X�m�d>׬�AV�[� �^�^Gx?ʮ������ø<�N��I�]�*w�EeYC(���-H����S����z+E�4_�y�P�<��ۧ������P�t�K�������p�<��
s����*:L�R��7�jQk��G)}*)��kYr�}>izͅ��P��HF���i!�`�E[��C��)N�5�������i%0)ċ��q=�qL��B�ҝ�齌s�v��$��a;5ܾh
p���i����b�}�է�7v�������>F�-'�����_��_Y���B��m��s(NZв���X|վ?'�#!Kd�5��Z�3�\��]q����#qNw��>M?�v�6��M8��sf�X����9�T�4��l#Z[��\��o��L<�2��gb����H�	e]H���UZ��d|��:k��S�,�z|O��4b+3Á�$T9��&�~��o���W"s���T�����'�5��qde3v#e�!������䯸�nW�u������	�K{:�U��!�r��I����;&�ql]��]�hb�L��a.�ݮ/�����P��6�(}4�Q_ ��5��DE �ٺ�jL`�d:��B��* +���	:�Y�v�r�pj"���cX*���Y�	���`4}�_2��sz�:��m�w�4-�����m�z��Ӭa�Q:�3/��nl�{ş�ǋ���gi�򨕝_'%�{��u�y��8Jo�-o�n��% }�KG�FF<����x��T���wO{���D��5��W����>l*��!M�����kr6������{f3��H�����\�2b���� E������rH�Y�y	k�2�u���}���`�M2�"�|�S��5�^�����0��7zs�fݵˊ��7�9xx[��*)�.N&#�f�����Ki+��I<W��g����3Fk�+�x�b��1�S!��*�6�
�t�@��@Ð����,���;r�ج�C0u�츄 8a]�ɬ~\+ݩY�����B �����nҌa�PC/Ybr$�-;��9�F;j�eq[�7��1�<���AߵQ���X{���2�R�Y���9!"�*�0��i�頋� g'�����$�`���֖�%Q���̉J���s�Qf��t+Q�A�����k��W��5JV�ƽO\ȣψ����Ѳ�x6.&��fv�m���]g˝O�ϙ���Q,�+���I�(��d�ӟJ(�������}��'�VZ�u�f{��K���ɱ��)��J�B��P��pe5���:���@^���ɗG�;'���7:�Nt��������{���8f�ɒ����*-xW~{��lw�?B*i=�J�U��,�l�DYeO����[/:�`�y�k�-M��wll��dۭ�����J��I���44�Nߌ�7�c�D�(;�_����G!\@-��a$�ßĸ���Ĉ�<��-��q���_�̓��,MH�P0��eׯ�Փ��Vh���A���e���4:xU������&I�,L%!�)O��|�k_�c0�y�*<t�/���囖�)���=O���,��ϐ�5Kɕ���5[���$�Z����'�snh�ȱd�l��B��^��T.8�n~<�7���omG|�e6�
6UQPL'O
R�1�zM���3n��H�>�Ҕ�+9n�FaLuš�
₞e�X��B��&��	��vo�qv���Vm����ĭ��Ѡ��`y;��p��?P�^�[�b��PU�|b��Md.؈V:�h�.r��I׆�N�)�wv��4~�+_������{��}���G���<��*N�$QUC$ew�d�?��}N�-�U�u�͠���c:��B؁�>F�*���'�J��A�L:�>��@B}�;*F�(\�[�|�^{KhRI8�cE	$��d	5��Q�@�Gk�9�A����(V����fz���\�h�v�O�f`#X�e(��A���Ζ�2�������}�4�T��>!� ��Ry��NMc��tm.k�Ρ�f��z�t���C���w΍>9qv�*M�_�,-C�9[`f�2y����H���@���*�f$�c�e�1���>6ѝ!�{�O/��xL�#����B������2��"r��_���)I.��{�"�Ʒ�^و0i&��7ɖ�@^M�`�~#��v�i
�^$�s%�`����5�D�; ����GG�PH�Gkq,��M�U�][2mr>��}��v�{^��� ݜ�8��Y��*SĠ	�$Z3�IH}|�5�@�U��������ũv#��wHCR������b.���z؎͡M��ĲC�c_A����`���b�	�)a�0t��s�����Tz�}4�QY��w���k���)�y��L�r��p�7\A䟦��3_Qw��È��z{�3�	ݽq��)H�H����H�V�k_Ϻ5�ј2ϩ���[c�;A�H��S-��|Y!d�3�rǚ�7QXZ��ϫ����)C��͏+3	��R�)q�"M�C+EJ���Yݙ
A"V�YW;�|/p 7�M�D�q������,���u�� A�`��M[��pI%;�Vc���Hu���ӅZ��v1�`/?g;\��a��~3��	Fa��o��/��  ���������5�����W��Ag��avw��Q�St�� #i |�]L`�"�KУ߫U06���$D%Y�}�Ma`�h�r��ע��NTW<��S׮؈d�ʬ�OJ�⅏�'�V�G#�_�D�Kr�N�����i��U�}�fؖ������vw�S�<-7�Z.�\�'��)�ܲt��Fa�c�/P�tV�i��@|n��%�y8����w/6��Hn�����s�X3���jaXK�ͱJ��I��y�s���i�Y��|�,��ofhW��� �h׭�=�&��!.��'�s%=D�w[��<���7�f��J֧�h�+��n65�>� 傴�\��
�kM�ȶ�4Bp��,,#�4 *
���4*tk1m?��,������d6\P4�A�9ӫ�rͥ�pD��[��69}���{��Wn��p���x�~(I����`3c�c�Uw��.� �Q��M��c.�{��⃿�-�`�c�"��=��H)��X ��B�5�p=��4|��6W�{K��0��W*�M&c��T��Dǫ��4<)pM]�ר\�W٘[ŧ��;�����ːs�6�#��%�Ď�����m��_�'�lxtl�Jk��	�ѽ6��n�ǫ%ļ�5?� ��ڛ��J��U�z��d�w�e�բ|��f�5Y���B�>;Ԕ��RDC"! ��mF,K�Et�o݄�qz�éO������Y{&
�-�n��]��=��*�7W�a?�b��ɧ��A�Q�7�*R�9-�ѕ,�ɦ�
vo�!����	 "�P�ɤDf��.��E����4bUft������V�9����?��p��2�� C�ت7���Zg�Vj�,���N��.���2ڇ�#���8�������d7"P�ͦy4���1A+���Xy�_6��x{tKUo6����3=��;���>�h
 �d��qefQ�աFU�̂�YjY���P� ɭ]�-�M��o�-��@�����wv�A��bI�@����Ħ.�?b;�_�<6�9��s��Ný�����A������9?�M�=1CL?��;L��<�QMnwzw��4`����LK1ؔPЍ�<5{2<�I�_�����z<�g������~5��nBK���ڽT�;�J�qX9�O��6
n�OCcnU]I�6����/I���}��[#��}���3�)!���h��1^@.t~����K���g$�
ևe�+�<�+\��������	B;:6,^�������V�)>�be���*����u�iq�K~��,9a��/��>��BީУ�T�IX�@;�QSh?���B�2�"~9p�4���%AU�>q��l�D�	H;����bB�&���c���昰���ia"�D&Z��=��}N��:!!<�4��ҝ�7����o	=�H��t�)��5�M��ӻA�F���T�zՌq���h�ϛb��=l�l���*��p��ɻ����Vׁ�����]�p��Z�ߛH$�GE���W�7ai��'�C տ6��t�չk���u@��7�0�moz�M����q���W�AׂE$�h��9o�e)�| Z+�r��ZJ��T��i��Z� �Ry؊E��� ��Ie	�3�}�� �f�8�!�l?Z7Y��e��,(�Ejp7(�n���m�]X�҇k�d��M/�WT	�Gt�)�F5z�_u��&XlxVHYEB    88c9     8f0���'��p(T�g�����r�,_��߿��d�O�����V�9fmλ��ƽ1Tw�3s04�}dz1;���?�v�HV�!��@q�65B�z*�9z��S��J��v\,��
��N�H�A���%"��|��iZ����E��Y�2���Ty&O��OjiIؓ�-v��+�Č^��:b�OYoa	�Mͥ(yߪ�ѝT�귝jcwf\����u^���PK�l*�N��{��-����M��i��1H�Δ���Ʊ��:y��`R�t��^�2i�����
sĖ����MbUQ6��
|?n�F�
@��h�.a���)��b������)F,F$��������
d��w����kaƹYB��4g�Oa*�/� �/���9�
�w�ŶN^�χE,���{g��{_n+����s'T�&1���Zz ZY�}6-g���S�7/ �%�|\p@��zy���#�E�l����FZխe�[�j�����߃�!�C��HVX��`�-b]H�Mv�m)y������8r]�_�o����v:to�L,qD1eo�5�Ԭ�����j׾'�=C�C�҅ߙ�J��s>#U��,��r���e!2�֗u�[���L�7*�.&�k�
�a�#��G�ksiU��u�{*�&10q�{� �1\+h1T�fF���Q	Fkd-%����b���xH_aN��5�T���T�����*����n�ݕ��h{F`�a�#e�`1���8���Tv#>��I�>�^��ӥ���γ�s�(Ӓ��zP��5��Y�ZM�%m�}�,=^�s:�^D�'�@>W��5�׏��O�>�{��Ъ�c�g�`�~J������B�N3�|�F$��P?�1�D�bd��vQW�����H���;�=�<�����|�Y$W)�6Օ�V�ho�d�ؘ�DZ��� �D";�)�oPq�K�ޣƋ`�:ꊀ�9�����:�!��c翵��k��9z�I�j5C2��`F�[T�P|�t�P�ŉR	��d�2��c[��Q5�.ra
��V��`�9�4�u�m���@s�O�f����=�0�"��ّ��9��tw�Z�|W��e�q��IU%���=���	�2�l�� W� |l݌�gb�kצ���V{�ל6T�9D�[�kj�����Vn&��ޅ�[A���n�t�������@h������t�f��'��[��MZ^���Y�AG��,����$�閄�  P�Ǟ��8	���<
3OJ&i	�j��t��N-��F��������{�-9a��������s-���{i=X��H�u���`���N��!跊�Z����W��I,�_��d�-7P�#��Z"& ��u���[��Y2r4��O�Ė�V��7q����V�h��` �H5��NHgD�,P�D�>{{�0��!����hY�d3��������lP�4�e�1E�.&lOeb`��[�@��_iue4/WOmc_<d"�9xS}�3�qI�X.S���d0��?1>�$�����X޿ŎB d�X,D5&P�����WП���3�_}�A���*�J֠�� ���Y]STW`�y���������ȝ���8{�JMP��ѻόj�ȏyj�K�N_Ut�5�]y5q����٬�����a�v>� �N�?d�W`�d��eU����@�t�e7�L�����I⦡�67�4�h t弥�ϙ���b�r(���L@�c&I� fB��BV{>��cC�� �֝���Df("������\�K;;a�C�~�� �J�'	K��q+~:n�p^­�P�v��'�]t���#�j�U�mٰ�z��_��`7t�\r��� V��boo����_GtI���
 �|wOs��B����O��6Gu'�]~E��ǩ1�@n��,���g�cܑ�E2r�h�(;�f�[b�R��K�b�h�#�{���T�}���wЂ��@�A�>�eg����8��q%�)p}��N�F`�Q�E֔*��ht���ےϜ���V�`��Ȝ��_����`����:�)D�r�[�h�?2ū��F��(,8�Nҁ鉌
,BI����D��K�%o�*�:,�b=��h�CV����>����}�%�zw%�AϺ�!�����ܘ��ְ���VC��<�-� s�- �?ȝ�����$����2�L�K�����ξ�'�qB�i����7���։���+�.JNψ�`4���W�]%�>��v27�