LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MB IS
PORT (
	fpga_0_LEDs_8Bit_GPIO_IO_pin : INOUT STD_LOGIC_VECTOR(0 TO 7);
	fpga_0_LEDs_Positions_GPIO_IO_pin : INOUT STD_LOGIC_VECTOR(0 TO 4);
	fpga_0_Push_Buttons_5Bit_GPIO_IO_pin : INOUT STD_LOGIC_VECTOR(0 TO 4);
	fpga_0_DDR2_SDRAM_DDR2_Clk_pin : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
	fpga_0_DDR2_SDRAM_DDR2_Clk_n_pin : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
	fpga_0_DDR2_SDRAM_DDR2_CE_pin : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
	fpga_0_DDR2_SDRAM_DDR2_CS_n_pin : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
	fpga_0_DDR2_SDRAM_DDR2_ODT_pin : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
	fpga_0_DDR2_SDRAM_DDR2_RAS_n_pin : OUT STD_LOGIC;
	fpga_0_DDR2_SDRAM_DDR2_CAS_n_pin : OUT STD_LOGIC;
	fpga_0_DDR2_SDRAM_DDR2_WE_n_pin : OUT STD_LOGIC;
	fpga_0_DDR2_SDRAM_DDR2_BankAddr_pin : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
	fpga_0_DDR2_SDRAM_DDR2_Addr_pin : OUT STD_LOGIC_VECTOR(12 DOWNTO 0);
	fpga_0_DDR2_SDRAM_DDR2_DQ_pin : INOUT STD_LOGIC_VECTOR(63 DOWNTO 0);
	fpga_0_DDR2_SDRAM_DDR2_DM_pin : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	fpga_0_DDR2_SDRAM_DDR2_DQS_pin : INOUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	fpga_0_DDR2_SDRAM_DDR2_DQS_n_pin : INOUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	fpga_0_clk_1_sys_clk_pin : IN STD_LOGIC;
	fpga_0_rst_1_sys_rst_pin : IN STD_LOGIC
	);
END MB;

ARCHITECTURE STRUCTURE OF MB IS

BEGIN
END ARCHITECTURE STRUCTURE;
