XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���t�R>��Wo�o.�_)̹4	�p;��*(�?W5��軁�WYp�|�x-����wP}'�}������q6�V1���	����s@�����Fˑ&X7��>^�eمG����X�;��Z0��ne�Ӆ�'�6� ��.��R<MalS�=H)�Kx�7d�D�� �XJ�"��ᷣD��|N���6Pˡ��Y���%�(���X��;����v{W��,�=E}�4�w{�	�8�sw��]A���B���rj�J7���+���x���=lk���[`��F�D`�Vk�D�j��C3���>{��g�p�ɭb�|��7����inA�v�C7uP�{J9���Y��";����Cgf���T:zÁ�NS"�_��b��	�cj?�=Y6���Y�jyc��2�(Cge����ϱﰏ��2O�����<�b�8ʐk�뜖�����W��,�l�"zM>��s��e��B�\�k��T�Z�3��(1{���W�f��'��̝�_���w��	�?��
c�Ԫ�&�=��mV4� K�p��{���ⱐ�	e�f'?(!���8@�e"�L��vvs�@?*Ͽլd�w�d���y��kȢ�t������>A�#�w¿wp������_y\NL��v��>`w��a����ק��ng��Eb"��n=Y�(�ZR$_o��F�B�էfh��9�'���4k����)�V��1��_k����e�HD�����ی�dJ�&�#݉][�3^9l�@kXlxVHYEB    4f43     f90�r���)����	q��6wr�@kB�z��m��H�:�n� ج���P�6�Uw��ۭ�g�)^*{L�jX3f�A����*^��ʋm�.]/R�#����ELB/o(�R�H>CA�"��cT����?�>���Xt�� �HjL� �!�u��={ ��|+ƅ���2U޹Z��ɘ	W�d/G�(�5��.g�Q�!������^wl��bqk���N�Ӷ/��	�[!�6��!�I<�g�~	r��?�H��!O`�f���)��> �0�%�F��IV�!|�&�.�Þ��ۻۃ���fw���TUn�X4,=.K~X@H
M	�3ϭ��n0��kb�R�)����Ԏ�r�@-D�z-�L��Z-��k�o��r�$�y=ӝ�~�9��e�6��������/4�r�ϑAWvkX	�<+�hd2�+�2¦�ˋ�E s�1�s�@������0�`��ˌb]����
JN%W�6Q�7��Qf!ޓ�S�~��!��� �r������G[�"wF!_��E榁�����mC���.�ڡ�#[M�D"f�����D{i3w�<����WV(��"c�j�*5��䖦{~�_'e��a繨}K3|W�ycA�5��+�.zS�6zi���>���P�|���!�*E���@]�<8�<�ӷѫN��cFj�+�ʾe*~�vg�D6UQ�[*�Qt'~�
=v"ߪ�������N N=
^2�����i��Τ�nl����o��6h���PB"��<c���LJ<�s8��>��U5��H�p��o�P���Zl�h3�T������1����	����y�\	�%�������Q�d�uӁ�K�8Q���_������	6?�!��I`�����y>עiM�N�F���"���R�x�N����| ����W���3H�g�ͩ�������#`���bU�ͥ9�j�V��/4;����a�����E
��m�e�Q2@8:�W[�`a�r��Ot�~����'6\Dc��nބ]��an�5%�u3	�'���N�`��L�j@��
[�'o��+�����,�s�l/pq��h��z��r
p�R1��Dd86�aj�Z�@V�dŗX)`�"e]�pŴtM9@J�o��B]����+�k���?^�h"�,�j��/�a��K�L��P�.�3+�}�UC	A�uؔVȽ唊t�RD��v�*z��U��&�K��cڛ�c��U�>�Y�M\ǅ��TF�k���s
��`�9.�]�%W�4?���(���%3ﭠ�f�E 0��k̋�Y���Uĸ߬�E���w�;|2sqо0��iF^��!���z$VN�?�4�8r]*H���٭+��@��ߜ���ܫ��P��x���x��t~l�LX	e0�2�����U�?��wem�t��FP�
#�������+��, ��_���T�D�UT�@F3�ؑƒ���,[�N���۩���`�L�_��z2���^ՙ�a�
y�6h%���k��òHsv��b��]����ɹ�XZz�8�g����{����VQ����,?^c��^5���{�<V��zU!��+6o��������4��I��A*�U�5�ڒ�$u���_�[}6����)|ٰ9a\Z��Xg_8���-�*����#2<�#�� ��:h����S��1c�����H���g�uP�h#0�p��ܿhjQˊ�����c�2���J�Q\�ܡ��Z(��9&=ۂq��x;�־̄:�%�{c��#*�*.�|�aR�l�J��r�p�n/�S�u^��vu�+X�DnLحp�����������c�&�1��O��!���X>�\�E�68��g���'����yB���J��S��B#�!��g|�[���q���< T�U�ΐ��*��c�_�n��`��$��iIX%���ԛdc�N��M|�+����z�Ҙ���6�s�М"��4p̈NR~�M��y`�H=1��y2����Ա!������y�?`/����$F8rjDlA��7�i��c�dKV��=��֯h���a\w$^�s��/=�'���e������0j��u!cQ�ܴ��|��c��y���EM��� yR���g�w���Y��cq��!/Ou}[��rMyf�e�O��؊6*.(�̅��1�ϚhC�cs����VW���W������W67����~��n;1�FpF'?���{�q�*�	���%�g/��XK;�Ɩ^Ԅ{i�,����φ97$����w�կ=�z�ū�8���/oDs�*4X&Dk,����<�壭 �|���'�Y���]�{�q|3*sQ�Ŷ�m���^���XD|�P̚6���Q��Y������>��I�g��"�*�p�K��EU��~썺��p�+�.�jK��7jd�l�7���-BYR�gt|��\3$��7�h��X֓4Bq0��7{
=��
�bIӑ�b&���s��Bֵ$V�ي�v��J��Br�#m��,��W��J_o4����v�,�v� 5�L+;�rvHs���HFɶ p�lmZ���+CG7pķ��x���۩�܎'��8��S!��l!���k����A�e@8�-|�=���/�����t��lҚo�8N=���f�a�O<lY�������>]u�i�h@;4�+���}l��I[o/U��M��If�=@|��v��|л��rԪ���EK:�~��H�S<�N�۷��=xl^B,Ȼ�r=*vZ����;ځr5e��02P0QxQ�Ӎ��		I�oV3*��`�P�Z�o���z�`u���[RGU�:$,�g4B쐏I�g�ytd��L���CL)Z�M�������.В�!!��|�K���Ƽ�@�5���Rϧ��ϟ��A�������X��.�ϲ8�m����4R\��͝�[>��p⢶$4dl-(�~3�����O��iȔ�tZf��c�{���?��i�4�v�[�T� ������{J���
%]jeEe�lPQ�qO�����6�]bB�ud�ϡ���e�BΏ.$%�����x���9|����.��v�����nI4�ӍA0�c=�i+v���[�I����v�����l"�;��X��Q�4�od#MLv娛�E���IqA��Ͻ��^�MK�R� 	O�Q�9����f��;yB�|�����F�n�JJ��ͮ��"E!p�p�%9[d�e}mƳ� ܵ*��F�<���`P#P�>}�������xD�~�����E���TⅨV��='�۸}��+ ��c�r��ez4Y�B����^͐ F�H ���H�,�²a�u��￟�j��Ѷ;ymF+����зZ+�ƽF46.Ϊ��HH7}�h@ű�ThY�y'�z�aA)�dbpc����[h�7���y��J���0
� �ב�C��6�.�J>C�v]�����|��'�~ơ�O�	��%y� �Q�0`E�t&f�T�cŸҮ��1a� H�9��O
hB��0Wj�4�C괋�N��d��H������a=4$nđZ:��!����(�<�� ~0Z�L�ea�HΊ�HC5���0K����b��-I]L���h�?%��33�� �=1����>�:6q)����{�_ƌ1��h_#�WH�;.�#M�q��}��)@z�J���#=�;e�r�C�o����G�@O;w�/�UW�(�&G�5�����|�)��\���۟2�z��>�4iZR'���� �%ЂX+SȔ�FY��p�a���^f�]A!�W��-!X�36�My�@!?Az���1�I���sA��ֱ��#��8��fgE��X��h�Y�O�$���s]j�p�m���r��4�q�����Y#�	zDCμ9)_#|~�?-ׅ'v垟�i���YM����N3ۗ���͘~@[��6r ��