XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��h@j������7p�<oL�yYs����#��y�5&�5mc���x^�V�Rñ�OCq+���L�� Δ�TA��-�XE�����<�g��e�]KM
m�j����C#�ԩ�#�����T�_)N'wj�!]���A��D
����µ[61͏���K�d�b��20S����6���q�R����͞��!��!�~.��(���G��'����N��j�|Cb#`�֔������"/�W�0.�n3��'De�t�:����b߄�59�!�}��s�ܒ��мv6�;+U�Y���>����d�LR�Ļ�՝W���@��"ө��N_Q�
�֫�}��]�n�ӓe�o�.��n	׌��;�N�ա��抬���E/g�}��M��7�z�����L�z�>%����	��`�	w$�Q�đ"��]�
I���K��J�u�~V���M��G>4�i�7c�d=΅D����+�D�Q�1�Ɨ��:=c����8_ù'�6�'J��,q���*�k�l�R�Zb���l�z���<��F��*o	��	��Ħ�at_��wyO�{Va�WZ����y���S�n����/j��6����Qi$������OUE��	���?�v��q6�g�3�������cg{}�W+1}=LZ'�g���o"����ގv�ϒQ*��()3��BȰ��"m�Bd"�͎�@Jy�'`/HޯB�I����v�3�W��<�W���}�t����p���h��~�N� �+@�"9�c��XlxVHYEB    20a9     a60U�βk!Pi^����>���
������U�x�WmMf�tV�о���%��Yb'�>zL\�dm5��)�i��,�O-��CM 	1��
��A*#M��n���I0x�y����˞	�4�����sI�:��g�bì�>��-��/��w�_�	T�B�z]ھ@T[p���˲︱x���4��1����C��BL���]M9yS�~����c�R���4����*���!۩2.�oc��H�wD_���J>�E��A�!|$8��[J�S��^U�����9�Vd����{nMPk�^ۚ����>~�o/jE^d�\��b5�cI�(�ɻIJj�`���|��z����G\�����@!�>�|ǲgT�,4�^�؆�"/�M�5sX��"]��ߴB�?�p-�$�i#6���N,=u����;��&�Ԫn\�������`�3J<1�TѮ��}?FH�ǲ�+-'������i�=�i5$3�R��w�˚O~xS��g���wQ��;=�<ꈨ��i�r.D���'��D�s>x��a�)�Ma#@|��`�B�i�:�w�	�g:P�	�'A�W@3�����<��i�dF��5U�k	z����oحʹ/vF��_zt˫GR����sXU�.�,T��Ch'���#���AJʀ�C��/[�D(�� b�u<�Q���,V[gI�1)n�@�I q��(�+�q�x��~�1%�w;�tȜ)����Xh�i�6d��D��r��)n�K������""�3?Qm��o���5��Y��-��C�`�5���/���韔J���!/�]y�^�Shb$�IW:�Ϊ�AQ���I4���.�L=1�6��Q�D�q$�ZG���1jO�����~Ӏ
5��h����K*M�	Oc)=��[=HCO��<ɞ|5�h�0�_�r[��ك8��`��� �^h���;��lg�������:o��ڽs���}�P�NM#tv�����o0���&ʠ�
o�[����_P��n�f��3�'���p���\���
@J�/�ܨYK	:��fIRJ�'�O.�t=�=��'�X
��¡eF6��z�ً�]d��9��n��ĺ!��_5�?j��Ԛeʣ%JLx<ԝE2���ϓS�al|.rm��oѸhAЈ���ڌ�@a�sKtl����r�y�N L�qo�E*�+8���g��cX����p3�îF�V7R��YsF����{mm� k՞�A�6�aܤk�/�Y]�i;�W��=������D�\�9��s����,:I�ʻb������#��]G�_�I�V�P�^��+dJ�S]G�eg��`���̹x����Z��������#��@̩��f��K@ b����H��OM6"#M~ ��H��W��w�Nm�ppÜ/E��3�A��U
���N	J������I\Z�������<����_���f����Ady�Ҥ�B����n�>cr��T�H��	7O��9d�FF��caNPzB�kӾm?~����G��عuL����}�sqw��E����p���~���Pu����u��W�^NV���Ғ���F�5�4"�Z^��M'��l��+�L�ă���$~[���2*6K�?���bFP6y��y��d�f�.�	fd����/���<�Ik\3�)k!�^�	������� 4����ŠjB�_ v�{~uMxr��?�j���W��G��U���U?�����V�K/C��&�5�	�����t����҄G#�n��@C�*]!Z"�C�Q�w�}*��	Fs�3�.�I���i:a�ko���0�XݹD��}���ź�q&s��M�0��Հɯ�	�55�v��G�oT�Ͼ>b���++.���X{zVMF�!��*!:f�������|q�y��2=��AR�aP�5��<S7�����c���F�^W/��?���3ʾ����̥�y�ŷ��x&ߗm,��b͟��XӶ�,�4��o��hͦW\��5}�yV,F
�Z��h$]o�%%�eb�r��t>,�A�0��x�+����ބcb�p�<�l'��&ϡ��׾��Z�] ���_�nQl��vδL{p���y�����Y#^����AoJ�QI�.6�`�]�+��d4�P��v۱�c�@���W�ć �����S@����^fl2"�#��)�~$)�ٳ�?�TMI�YLS;�L��ld�qՇ=��r�L?2����H}�>���L��X�ou{E1_J�@�Y�0ۧ�l��z@[�f��NU ��j��M�ݻ_wL�ҥP�]w8hriIx��J�'˪��>���&}(�8Lm/�N{걡��WtG؀��H-��6�`�3IQ������lw��確R��OF��`cs�C��J@+	]\�?�����z+�C�\��Ҳ�-�C�6�
#h�<�J˼6������<������U%�xbj���`|^c�W��("q�8���}�<r�o��!{�����A):e�:��-�����z ?n@�m�xE�(��a�KO"({{�В�aށ2|f�)�&���v��8��ZqViX*E��,SuO�{�A�������S�v�4	�ް��?x��ȁq1*�����S�����#i�