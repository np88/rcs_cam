XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���������ߐ�D[���?$�jϿ�RR�kb�����Ͼ=����تTd5�n?f{�R"P��p�4��h����������oHn���6A�&#�OO�H@�
#xlx���)A{�SOA��K��F߰	H?���/�iȵ�o�Gyz���<�<!�=��b�r4Jp>>aq�<���e��H�#�]�����qI�$0֑
�Y�~����cy�j�fX=�KK�ĳ>���d�$��b=�O�����5l��`GH ��d��N>V�dj�wM ��U>Jkl���β�6ȡ�S:��(���N04ш����� X�P��T^Z�x�	��V���i%�����0qN���NJ^ C��W$�����K"ǧDE@�d��߬���9�؀V�d�J���sZ����R���Rs!���je���1{ -�%���Qﰼ��Z�.��m�ç����1ؤ1ۛ�ߊkj�<W�i"��Cǳ�r��h�5W���0X�3Ȗ��J�l����Ĝ�H��0%HQ3�\����	jR:�]�sM��Žyhɑ���m��)xLZ{$�*��|&3���6�Xf\��W��@F��M{��ol�<�"<f.�3���@�=��g���F��>�l��^A�� �)�ڍuO͏�{:Vǔ�I��<1�UJ�\�@8`<E�PZC�<4k�j�l(��h�_R��\�)�a�}Kh�٦����ǃ�W�R@y=RJ���η�͎u7l^j 7|��N��~txA�b��PL��PsuXlxVHYEB    1802     830Y65�[i�~�%s��Ӆx����~�)�T�>�;7���F0�:���Y�[�_�+%Mk����]�Ǆݗ�l����A�&���`�����qȆg�G�
GOYߙ�����QA�����
	 i �4�|Hjb�{�}��>���C$ w<�.b�ԳC(@�9��ae���.܃4�6?/�/�-�N�]��"�) 1�\>�V�L�#_*TfH��Idp���4ዦ6�"l��;�?|����#q������zz�V�s�YHt���w+H|�
"hy�w�k�.��p���;���O��.s��KT�����*X
�T9!�s�?Q���C��5����Ϡlǅ<��W6�_�X|IZ�b��iY��S.MB�^`<V[1�X�C�
ސ�:��A�(�
%�qa�g���u�ד
@0N!([�G���j낒�x����ځ�%I4{����!�_���\ǹ�Q0z�2��FaK��U�͛��TH-����^:�m��!pP�=�@�{�hՓ/�Qa�ڶGt!��h�ү�:�t�N�yH�bR��%��fP;,�y)����D+C�.����$+���僟���~'�(�I���O�����������r)ᇫ�{�(����I� \h�1�Vݕz[�N��M��G�4��-0(��"���)�v�=zL�E����Ц��Vף�M��&ň%�Ɏ�^p�x/Ը�?���"�D��8L+Ǿ�q_{h�3��X���� ��`&��A�v��ف�����G%8��ni�E��<GP�kIB��\�p#��G�G��b�K�ٻj�L�6	��� =��P��s�h�9e\�����BMF �f-`��A!����)�#�Y����)����涔����8��Fr����`�*"�-B�c��!+?���8��#�;���o~2�k����Fu������M��mLA�; ���7���E�kvo����Ag�p�L>��l������
�����f���9+6�gW�\��IA�xһ��K9h����,�k��Oh�_m�)ޑ8��EP��炨�.�n���CX��n<��@���mؓ=��Z��Mȼ��"MnD�&^���P]x�P{:�h,���t�b��_�������H��[�$��w *448��Z��S[�H$:Gh�&r\����I��v��ڷt<�U�c%n3Y�(ӝMG�=|1
�s�.Η�NZ�%e-��[_���:����\-M�Q��ys:6�]�,��$1P
��e���i�A��o☜�#��l�P��S��T�m��XL<�o�*��D��G:�9�y�Ck4 �R]X��4�%�M&u�S�
ɔ�b���D���QۖRj#(�8�ȶ�&��\;m4V	��ܔ��0na���������^,����_q�m��6�8Tcd���_N�ްO�����}�{W?N,��˭�\�
��_&��-J,[)�5��C���W�V'h楶��~��NR~o�k3�`��	�B�#�����t
���g0��h,u{����d 8iRM/�#��6Z�Q~�A�0�=�?��n�cx�������Y}rؓ
�e�"��v����P����s8�>���t��#7�i��,'��U=����Ow&���G��{S����-�^|9�'N��^B��3=_e��&p�F�.���+"�:�~�h
O���H�w�[�����1������YBJEݮ��aZ��@�V��Lm��Z�d򤣈�>��y�^��(k�$�G4xoX5�u?�JoD�� ��u�#��ߡ��u7�7��>u��"S�w��0q�թ�Zi��>b�e�����1�)U�~���_�@��#?A����3�����\)~Y�Z�<\a��b<P�Ž.s����{r��Ui��J�}6p��_	p�e�-ݜ���w��}�[�J0���j��v�BM
���㩕��T��pd_(l�Y��䝡�AY�]�~�I{��� @8a�'��gw��u	H)�U���<"�3�"����S����M�>��l��Խ�<�L��� pdT&��G��~�+a�