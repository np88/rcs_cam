XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����Qd)��eUο`����l������VN ��^�5�a�:{���^X w.0�
Ue���5�<��^V\���OG�jT�Y�	�f!o���y%Z:�����r��=���H�^Vm��a�i�����@��o��~�Es'���E�?��������/Z�4�9*Aw���nQ��y�M��%�0������Qly�aſ[�^��z�����@�ؼ�!�PcB�8ؕ�8޷�Ot�vKS��ف��C�)�d.ޒ`�}����w�Hn�K�9���n�t�X�5���oE�+o57� ��U�A�6�%G�M5ʀ�N�'hM-�
=�ͮ�� Q+3��c��'�-Jq�:%o3��݀�ti�ci�h���fA$��iъ4#���|��-\d�?�T�qV�#�`���Y}g.�U��>{�M�M�0�Hm L?��~� �\�&tA�ay^~mX��l�z���B�%y<�a��}�}�䨉E[�,�P��m�QH>��������y���}]�CH�����P�cH��.��ʭ�4u��{yz�i3^i=��q�b�ie�;&�"�S�h<H 	!L;[?د9�4�2\���Z	���#g%��u�Z�?�[���Ww���_͕G
"����|i�
�;����x��'v�YPM΢}����������)Y"Va��駹=��FŞ�~��aM9!}�Fl�
X�Iz�L+��_i���M�~o�թnm����
ry+[�
Y_�x_>	�d��+A��茜��A�%�M�XlxVHYEB    fa00    2030�kf�f@&�2J�����Э4�Q��ɣ�r5�G��A90����d:r��Q���*J�2�qI�AlZqX�hJ,<@�Wìcʟ�� 4T.r�����%r��|�{p�!T��?����[� �3�)�w���=��eJ[@e��`�@;�M��wBgy�/�-��iķ�2W]�2�4B�ʉ�l.�{��z{�z#X���������q���n�ˣ�.�yp�Z�yp^ZYU��!�%u���lk�i�tw���O���0�s�,b�+%��gF��?FC�l�ܶkD�nF>�[]�r兊�]/zkV�A;�}v��F?*�Ã��/M�Q��0R'��Ū���o��6�N�a��Elql��$�p�m����[��Q���Ow��Sk�V��Z�H2�mg)�r�<'�<H8 ��eѰ�����=��s�m��ƥ���i��������`g�=��$�,S�`��.����$?��L��n�L8��ZY�c�ˑn�x���x�4!'��}��#�[[��9�o�b&І�ldE�+м��~Җ��M�4�A26�i�	G�U�@.��N��UKǍ;{��uŻ��j"2گa��H����A����p`��L�nN�t��igѬ4����ZC\�K�}ޠ4���X�i�.M�m1!*܋ஞ�&#�&��XF�/"!���l��uX���=H��f+��o4ƜfށN�>�v�v0M���H\�sW���A���{�Q�I�.�s��/p;�QS-���H�|p`��}��T�����ѫ���;���&�q	��o���T�d��Y�RR_��*�kzX$�G�Z�aI��2��~i���q�/�*'%srq���g�C.kju����50%29u����69����Î'q#b
[���wV	<^���Z6?����}���΃�g�6ǚz�XC1	����
�N���E�����/8ed�$3��Es��㧭ك�"t�}o��k\�������1�&���:�Ӛ�o� ��e�P�$�WU{��2$V8w� �9�.�W�/�B|��(�F�G.mNm�J��G�/��6 �쳓}¨׹���9�cF�D}���i�u�L�mʿ�ܭ�j�f+{
���s�'8*�j)`�@Zk���mEqW|?J�n��9��&�iPhI���O��c��`��P�X{gYx�m#�����3 �$4��$��z���	�Q��'Y��d���>�i�c`�����������񛤩�o�&ځ�.�ԭZ��mG���4���@�0�����~�~l�h�s���g��|d��M������t���@�9�1
qr
T��w����)�p�B�'`--���I�<���I�s��4�r����DA�~6�g�$:�o���b7����;k]�N��|�>��Y�V~�7��'�z#�^+���E�Fd��rѼ�eo]b�OQ���-z�+t�D�ʎ��]��?���o��� ��o�a ?�U~�p�@9�^���@��B\�l�P�p��0[�k4p?C!O��������h}��'��&;P؝K5�ay		Zځ���F���J;G���A�8i�&�B=_�i�,�}b/}�K}vn^�B����F��L�n]*f���� ;�<���FH��s+O�fݟ J� �W;��cR��f�u���tͲ�rg$�������5�`!P�Y�P�'z��i���������p%�U�p8�шABQ.����Nb�u��,e��$��5���	#�Dh}�D.�E����)=ŎK���}~E�<M/ɽ�D��|n�޽�d�g��2@K�r�X;J��%�����1~[�u���/j�Re�J.��v���՟S�W���N�u�f��ظ �=?5lӦ�#�tv�{����]�r��eG���ķ�$��p<�iݱ�(P�ٮ��� �P���:EUŸ����4y�6�Э	9@N
�Ad���������7�Б�����ml���cT"ʤ��/�5���ض`�����A�=�����S���l&��f�!�萖���h�"Hz��5WMa.A���uw��y�`�
�l���0�Pk����)�}B��u�\䍐���(�GIk�~��kա� ��(H�2�P���֘�)nr�w����r_�\v(��L �6Rr��{��E)p)Ƅ4!�OC�>�\Fϧz J.�!S����ߝwo�׸�ǚ�IP�X�h����9fo�1���H$��:�ܒ�b�#g}V9��y^���v��L�h�ڦ�GP^�h�T�v�����$(ߟi��,�G��Y,B�-݁�zD��|ԫ읈Y����!�����m���e	��F�WW\�LAW�j��R���I��)�h�v�x9�GF�(E�p;��ݫ Ń��B�r_��E����w���)��F��-^OzNc�<$fyak JDH��H�"�{���u�z�/�"#��֚;nJ�L)䇼���/K���vЮ���v�^&J�fvb�^0�Կ��۟~��>2NaѪ{�{����^u�����#�KխPÒ���dx���7���à��5���;��&$yBh}H�̢X����`�_���ҍ����l�Q�hW�����@��B掯|���A;	�$
I�<a:[s��E	+�beM�B;[���!q6GL�<�x�Am�E/���$�?"gZ���������.(���%���Z�'W�PkA+rF�hӋ��ם����j_�1ȝ?;zԀ�<�~�S���G����8MjS�f=�����)���U�_qyt���ĵKkl!�w�.n����L�ed_!Rr�i��GU�> 5�ł�!���u+�$���i%�,���}�ð�H�}-�H�/����0S�r!O���(�è�ʱ���t�s��{ivz28(�N��Y����4�:�֖�Tبl4էQUԆ5ؗB<A��m�3o"+�(A�tU=.i2پ�y� |���[�v+�r5; +{�"�pT�e�<��	��i��"�P<M��2Q��¸Cӥ�>5D[�����A��%!j��ѴqƘ|N�T�ˍ ���O�aD��a`b�K3�&�rU�%�r��oA���t�9h����t�Tr�a�ͷ,HF��T�e��fz�| �F��S��O_���=���J��^D�>g�F�0<�N}�Ej�0(���9nE���ng�r�`v9�5�Ӟ@��0�p����~Bx`�d�}rv���!�}�p����l<��ia�t	5���>"�`�rlg�
Kn
���|�I��`�E��/��S*��w1���7�mI]]K �)gZK���O�����jg�w�=Bc����|�Z�n8��B� &fzαK�Q��¯A���a�|~"��u+��	�.Hdw����ު *]V�3rA�_���ąQ�O����r�����?:�&]*%_���#Yǃ��f�Oq�Ѩ�T�Ε�m�K�.�sp���|�9�3Y�q�F�����ݝ�I��$@�Op�ځ �`/S���KB�3`	JT?���(<?/�����z%����3��;8;6�>�o*��mz��T�$�����Z� �td�{�c�W�zVk����5�
4�
Q�ji��) w�4���8��5`����V%��*XRl�Gؐ��{�D�ĵ�3B둀��C ֶݘ[��͒�����x�R%h4�#ܡ��jy\d�O�H_���g�fA8���
;�1O��۹0F~�u�R��,a�=�[��+o����AY���c�^j���xSEؾw`��*�8a���s�a�<vy\γ_��,݇�$ ���6��q�i�+�"I�+w��L�]�~^��O�K�c��Y��.��B���fXo/�8E�/�������)B�L�]�o��l�W����~f�~��S�n9� ��G��	D���V��>l�[�cC�o��e⎐O��#<Mu�ס�����T���1 �f��n�n�6��� /����x��f�m8����f�Y�2��=���w�|a&�ʻ �|�S <��aD��H�p�,�#�uOg��kC<��������|��~HI��ޗ�D+d��@!9�2un�U�S���v&��) >��5���n�u���|�W�㋆ñ*�M�3�>0&Ke�I7�sv�������Nr񀴉��ކ�N�ig=z�oZm������..����[��Kn�>���5+����>ŋ��>���zF�)��%� ���9[>Q"҃�c�t��t>5]�X�{�EHR��0g+�m�U� �/�! ��HBU8=V3JY��7^���"�Fw�����*)��+c(�{��v����f��C�t�hx�:��Fg.��w��=A�	�巜�����g�=�v��i��<e��
��q�Z��i��c�"�ϓ�m��/��_�}�;A�e��2͇$�9{�-���fZ+���_���qa�2�j�I�bn���2�$;=�!�+��J�DvJ��$: �f^=��(�����2..�)��P��:��d����[ ���`ʬjo>6tc���Q�<�_֠��0Λ@>!Gո��&e����t �6]U�I�q?�2EE�te�w�/ʑ6�Jp)�lȧVPP���J6���5�㪭��	4""8:܈�&@
&�J]�kZUWf��[k�)��Nh9Tq5}��yZ�vMچq�U�k6�'u�⇙���޳��؊�Y��q!$P��nx��k�Ȯ0�u�:hx��a�%\�J��vÖpN�W�s�����=�k��!��A^#Z�Ԯ�M���z�1��m*P�|��fCBRu��xs���ȶ�'d�T���IB��n���&��9����ѐ�u�'�d�r$����E��h�B̀��xII�Ԟ3O�H��R�/����_,�1��3Ѕw���m��2���#��۫0=�m�/;n;t]��Bf`k�N�����.eQ})�M����>V$�oړ���Ǘ���Ǟ�w�� �C�����@D�����X������E��?͹7��~�3~���-P�#O��!�nL���?�5��U�c87���$���#Ǝ�x
=S��a�z������Jg5c�\��]�XG�Ciڔip����E���nǾ�-��7��[�YO�>��'���e���[A�U�14'���<�5����O��3�:|MS�����`�-M��YٶSD������w���N-�� t�j�i{A��`��Ϡ�	- zcV��bo�?gA����Ij�F�H��{�dp�N8��S3�.fC�FZ��P�u�>�!���'�sm2��w�N���:�{/��]���~&�ɼ��F�O�4���*��~��G�D�*2Z�D�:SI#��Ѷ Qr���fO�zj[��Kf���f��$��U�4�`�Pi�¹�����푚�"�]�?�Ι����cBQ)M,�9�(�v�x�vЄǼ�թ�R~T"��;Ť�!`�YǦ�%0H(�(�'G��$A"�b�S�b[�,���|%d!�K�`�@���G>� s�
��p�5�5u
���AV�ד�V1��6F���ys��!�O���[�V���;���q �Ҵ%@7�5wՖE# e7˲$�p��tJ���lWIc��hDN�]R�_tEP�#�>$��`QƮ�N']\H�����לE�p=�{��Q��3��:%�!nN��VZ���b<��ϒ�F��ۦ�C���x�;�pw�jQL�\�����m����:s���O�D���Y'��h�
U��c8����v������q����d,3�P�x��(��3 ����@`LYjO��mez���rU2z�*B�=tA��o���lPs�[it"K�v�ا9�H�>|��u��6�.�I�֫=�=C{�-�gB0ꢅ���7�(L�������B�%/��\��c��]pևR��p�q~ſ@�S���HYYgN�Di�{�჏�V�z���7���<���Zc��-xn����=�$0Fo�N�>P�e�s#�g���G�Z6��~�햍<�Ԧ'��b�F&C�d�r�@�P�-Z�NB砼���`J��=͉�3S�Ҵ�7��S��B�0˱7���n�B�|Wo�<������V�I¦zt�):|��+�_ݨ�>�/eJF
��:���ld6.�",X�pXδ��������P^ф@��\�!��w���qI�����Z�x.K�V�-cu�d�S2��r�j���`�r ��T	}���e�y?��_3?W�%��J���Ɏ�(�={�ml����F���̧�?wuo:A�ֆz�c�����su�[�U��#�Xr�Z��?F3��!]�F�0[��z���E�`���a�4?��F<�{��qb��Zx�^�2�N��؛�����K@��:�Ć�ݼ�`o��`[Z|IuoN��Ek��:��ҽ����g����ȑ�F����=�+�jG�k�am����"v��ڔ#[����ߣ+��A�J5=�Xͯ�ؓJˮ�i[�����1���o����{ ��MBsX<��Xጮ4��~�rfȯ�3��~�p����i>�>/K)�?n�ې�#����0��sK��Cf�輋���UOb�ُ�dަ�Z�,v:L�?�ʼ<��7���H2���mP�3'Ĭ1��
�Ԗ���D��[HG[�bɘ��?,�G 4N�A�U�W�wp.i�����PwO�U_B{4�B�U�IM���PS�>���cP�o\uB8���.�Tj�3���㑠RE���Oڶ��!�kJ��:*�����V{�'(#]#�3��Z����A^U�ͭ���A�����������?���n���������y9�N=ltM��|^hR���V�fff8��g;�*������3-U���>���!aI�Xd���+�?i�}��?�:'�9/�	V�6f<-vxAf��-�?w��Փx�cr(1����7➧��ݿ��z�����9�����p�.�	��������~!���9*��{r���b�?�m#SeXa�L�yjm<�f�@P�M�Xt���8E\X?7��N��B�@Oo�����o�q:��B=��@��K9! ~�Cʷ^���U���䅉��FF�y�y����pLC�{`�e�
�|�����+�9�EP"C����ïo���ucm3�hr�qe;��ƈ�G��O�Q�����V����Khl!t����,YD���Tk&�"�}�'���ק9[���g�ت4P-3��G�,���%O�4ut�-��K�Ŭ>�nT]o���z_ֹ�r���V������#\�ς��@�Q}g�]_K�/X
Li������^Y#�p��A)��"4��`�T��Y��¡�m�Si�e�8����	�ÉWZCe��A�S{��ɻ���[9�@9�RfKO�rd�[��X���`ɨ���C2�,�x���Tmu��9o	��A���w?�?]�f��1{�A��(���T�2��Eu�im>��� DG�0�r����n�	�Tv�q*�Âp0�;j�Җ���Q�oY͐b��Ӑ����8�fʋ�������x[�
���y���:��SƜa�$-�Z��y�u�\h!����j�NQ,���=�1hT����%z��wN\p�R�ɧ����(�1N�������(�>�D�P�V�f{�%�F(6�eu�@��v�Ł��o����$��[�J�@Z!c#�6DiGU\x8Cx������� HgR��~ej��w�h��B�o8Ațר������oUf藺���o�ߢ�(�et������wn�U��ـi�w����Z�@�S�Z�YU��< M�{@u��{.�듏�:�bX�8��w�db&�b��z�֦|}���m$�톊&���Ĳ#���G����;4q<Ү�rG���`�ܟ�`�$����tM���$���W��F:����H�e��N�0��N��EV�xxA#.�S���d@g�0(K������1�~�M�cY��r"�W�����)�M��������v�KU�a��4�;�Xs�����k�n�6�مzV+R���`\���K4:�2`�����@�?w��`xq�8�XJ�`��6wCXIXlxVHYEB    9620     d70��W\/�*���,��u�[��e9��,s���i���8�"�����]����\(V�-> 4���H_��5��'��43����ۿrժ%�ݔVU����i����y\0v�^B�q���h$n����#''�ѯ��-�E�W��}��y-)H�t�v���o+-����HĽ��؀�0��Z�yzp������Sax��x��w��Z�aX�a�ڧ����\��$�O���������i�w��m+���k/���R����J%xaZ�������Y��g�jS�y�-_�k�z̓2Ȃ�
%�D��O ���3h��>�F%]�^Q4��%�Mx5.�Q�6��[Tj�ds��������q{���3�r06~��A��^�܀E~�C����y�Lg���	qy0D'B���s�.�4��5vU:�$w��V���O�+j4^� �ƣ�*���Զ�Z���Z��AYLQ���;Ny����uє�%��/c��-�ڏٓ:�Đ�����޿B��"b\o%����h���53)1>$Z��{j��ZL�>���+�gј\�E<���w@#�H�R�n;�j��������-�l�/>���bi�s��m�3t*AHBS�%��U������<���kq��N���T��l�1a�	�W༼�l:�CB��b�\���gۓ�� 7BLmd��=�I�;�d�Qjʁ!븝�i���lS����Y�Nv���
�G�.ΧZ����X8B��P��]scg��Q}�I�e�8`ǙRƛJ³��8�7�Vo�j���`8z��!I�PlS��o��Qg���y��[G��Q?��a���s�9\p.�M{�P�4$z��\�~���q�K����>�	^��z���O�v��{�o�8?b��*�:~n
xO	��/�u��b�soo��-D�II1i�M���^�*Is���ihKn;#����6��e�s^Rf1�rR�����2i���"�$#n��Z�g�E��?\H`�����hj��M�o#&�U�@�^'OO�ťP�`�D���%�~��Į7i(�ɣM�w>����2��)bVC����KiZ[��3�A,�/_�5�^�<����/������l�O*�	P&�E�}<�;����@#!� ���?�/�LI�K�vI�w��w8ݢ%�UpK� �<%����Q�����X���I4�Bɿ7�;n%�ĺ<�:7sp��W�c�x�z�=�vq�d�U5�T��qg�ƖG�у�e�^�yg
V��������T��&�%��H�O���c5+���0�`%�A�����!^4o�����"	Y�+�EE-�>��R�w���<���{}՚�}e��S�$��QV�\�8�o����6"Υc7!�
S.�t{�z^��
eG���$���'��<\)ӷ�jqQ�z�:�`��xp�h��X_�7�;ؘa��;&h��
�X�(ʊGt_�]�ֻ12�@[l�Xm.�x�v�v�m�2�j�$˄�V���L���!�
���.$�M�y���,�2�^��Y8U�Sc�9��3���i֝�.� h��Si���茒Si�S"}s���C�q*�˩���*(�DV�p�4{_2�=!+MB@�d��|I��Pd���xa��D��̀���eJĩ��gB�$o`����nz���V�O�	߫��]f��Ai4��\�X܈gy���̅�$���qxԉ�W���4�5<Kw�-jQZJ�7M3)04w�jj�>i��m�xf�i�y��YsĘ�ZV���7 -���Ъ �d�
t�t��o�Hc��J���n�9<�6�.Wȯ5�FI���Ɋx��j�C�b�I��C� �.���M��\~o攀�c���H>��Ysb���0[g@��.��-
)⭛�xǸ���o3n���U���x��f��6C� ��� �I���(��3����T�+����[v��>���}F�Ā��;ݝ(����,;�{>DT�9�;/� ��A�t��G���g4�4��g��g�E('BCk+FXo��`�@��Y���M�J����Ց����}�=ۮL��Z��P���>�ʼ#�f�u�������½�S���:S��Q�i9]0��K�%/Eܨ�q�U8�fٗДݾ�~]Q;N��U�� ��E�Ȳ��Y]������Oh)?�Q1�:{�x�z4��]myb{�\�6�*�����T�A1�L{���!y����54��_Y��r6��So�a��؆ǅ���O���/�#��Y.�H��JK�.�D8#����V�h����r�I=�+=8�|�'ga)��E�����Ʒ6��
?�?
2��ZЈ�ҵ����5��'�}MnZ>�y �MX�w��Щb� Ij�l:0�.�D7Lئ6,�ZU�	0��!���l�/�u�Z�j~k��Rt��=�@��e�\�*YR0�ݰ�Ht�8����(�"n�y���d�wt깤��	tw������@hFЇ��'��<���:�x=��s.�v��kw-M�("�Ny���/���%p�� �'F��V�U) ���.<rt+���P�y�#Y�k��z���eo�E3��&��qm��Q��4��٢�0$�an�|r$� nZ�R-�Y��<���S��ؕ	"Ǳ�Pƴ�ܴ1w��SZ�-�D#��z헙��i
��r.��t����B�i�d� �����iy@evs� 3�C%�m���g84y1��;��Gu��ȇ�n�c��h*���"�18�Qg�6՛K;���g(2!�kףi��9�84��q�b���Bb2�3�h�l2 J��o�׿D?t���tH��&կ������7���[�^3�&��y�É�3��8�t)-�ca�f��j2�)�(J͂�=����Բ.@X)%Z�gO�"�Ғ�p����u��4���wN��� T��p!���dBSuÞ�����54%���mbO!pc?TVhU�����֟�4�u�ڦ����luF�<�5G8X"��	W]����jc[,��]�^x�����x3�#K$%�T|��^���wL��JY��W��nn*b�d9����U _��_�ZR����A��������_*���.���n$3e�tԃ�;�۴kĐ��L���M���_x_�ǅ�����	r)v�6��~��8��H��KdA62��$~@�ޫo�)le�P~@Ed.`_�s�J�F��F�]	Bԅ0M���]|�#�`�������j�	޵����w+�l~X���	�@F�<�0�.��1[F7����j"r�?3a���Q9b���C��a�=�7+|Ro���P]�1ZY���i���vJWQ��	�QK������(�?̂%'&ЉN`t1F�!�'�5�����hX{Lߜ
��/_��û)����'8t