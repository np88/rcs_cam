XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����]9U
�	puN��(�ɂ{�GZ�z�oC��pV�y��K��Jm'Њ�6t�����f7=���l��BV�P��r��E|ؠ�`��.�q�`��ш1�`� /��Fo���;I}t"���S����`�����@Ľ.휭9���=7 |���
*X�2޵i�A_-%r�c��zf��tq�]�2�n� �1�S��h��8�*Â?��L�N=LA�/�W��r�'��~�g
Q/�4݄������ҵ���qߢf�.P=~ٌ��0Ԓ��8�Nh�S�qճ"z�U�� �)��-ߦQ��o�!5[b�^v
I�0�U����:���x�|J!l<K��s��� ���´Հa+�����i} m��f�9L�.�
�e��������Ѐ����f7es�~�x�	}�m�Z��'��)W0��>�d��|f�+����?w5Kc��9���*}�x�_� ���w��xA�D}�ob%��0��3֏>
����!�)�߁h��%�L�j��������V�x�|�@�kRꑲ��N^��|7N�vU�����ڵ^gŋζ1�s�lY\�;~K�kC_��V)*����fG���˻a�7$�A�_;\PB*��$Ps�OW=Ұo�A����3��˪��>�$u��7��Au�r���s�Y��w��L��u]Ə'�p�8��6zU1���;��Iܩ>Zp����^w-�P+���������O��{���e�X������Ћ�AB�LH	���XlxVHYEB    549f    1060��[fD�;��p?ݗ�xh�8��s,Oc��������3p^�n������6�jd�R�T[�X~�a#��r\>�A�&���13y-QS\��Pٝ�D�b)Z�R�\�,��B��B���e�o*�m�J�g��+�q#Z_��v5�f0-�>=t������kOR^b��u����w>$`��niҳ�E=�b3�^��섐�����W�Q9H���2@�G�	�68f[�콬�W�C�í��ї)k�t�A��"VAyTV��Cg�DC�S����ߴ\���Z}a$`r�M�͜��N��.㧯��Xh�.�/#��X�
��kͬu���0����w�H1հ�kf�;���
ht�$fMe��
z�����쁗�H*��!?�7���hL@�B�|�����Os�����^&T�X�%�C�(A�|���N��e��cq�J�n��M�s ��`յb�J#B�6�}��]�����)G,�ﴻ�(@fJ��oH�����/lK����V3�ꡤ#�ƠT�sk��2��z??�]ФjS0�#c�z��M��+�I5JW$Z����P����7��5�aE�t��o(��J
��b8^�ȿXC�A9�IY�Q�*m��m��Q�_'����︮�ƬxVta�]#��g
?ޠh=��� ^4{jn����6����9�|�B�9V읷������g�9��C���tB���3HIQ;��pjYi&DsǱ�N3�ʵs���6{��b��̆��lmȗ07�/x�.z�ٴ��ط�<�p+ؑ=1ʪS���<���U��
ᕾ��ۼ%�7�DxF�\��>�.O]d��׽w��NP16S��ZO7�{�"T/Kn�)w6=������t����l�ޙ�X/�v���A{����x0"o
�������k$_/k�wZ�9������i;�OH�]���j@��Y=�٫��{K���m`�U�Ej�'�V��u�.=�z�E�7�=uc%A����ZѮ����N�"�����%�a�i��ص�Z��ڭE`(���k0=e�'
��Cl)��(6�)���7�i�\�N��G*WA-�+4�6P{�_���4�p���t�_FD�_���hM�$�1�@!>����u�&�F�]N���5bMv������3����s�?ݞ��� ǦNd�}����]��|����#��u%�O��]FI�@0B�
~��	�����Rv���x�&�{�������U�v��:�X�#^�g���b<�7�ך�4�X�KEo�)����la,N�6f��ӿ!����ۏO�y�<L��+��3�$���v���t��j�9nxL4p�e�l��tSF3F"�$� ?�,��ED�	���
�YZw�C`�]p� PO2������h}�`�s	D|ӡ^��a�p��X���J
qٗ���e��zǸ��}%lG6`����67�g�=zC�wW~�"��5�\W���0M�]2�Sz�-�k�e�qR�:���ܸ%���4�'3~�	"�B'�=D$�5���>���"�aV�	�^��"Ic?=b��fAJP�����7Y��j^N��Ҏ�@�U����hhA�=�*k�Z��ƛ��Y[㌋�����7[
��>�Z�C�=
{}֭�(n��s�O	ɠ/�a���
����`iz���,�W�x�C�7�.���V��|�X��L�F~`�� "��XR��z-K/��I�`.�f{�!)}sA�g��Rj8�!G�m��oJ�[�y0@��3`=�#���W��j��3��ەG�e.�j�(�������qDF��އ�Agdvp ��T�D�lV�t{]~���P���}��w���y����%~wR+by_�i[�����}S-�Y� J�䨑�����Ϥ�T�r�f�F����!u��55�l8�4�~�)�q�rW�����[>W@�����V9՝���]����'C���*������"���f�u*lb����,�`��\�ͩ]�#���`���U�r�E�8��Yr�\��r�������Do��T�t�Vh�_ 0��GSwnf�=�c|�fC����0*2�+&#pt:^�5�N ���� '�H���oc��;��ٕ�I3���9t8<��4Y/ٕ�ŗ0Uj�17�m���i��L��Cc�` 
�I��@}j������a��
�Kkɕ��y��*�-4��i&oi1&���F��8���`�h���WR�H�p���&� 9��~j��=��O뗶ޟ?�JI�*�  �����`�h�7#Х��Y�!�#�p��'�x(�#�N�|�D\�����^7�wV����y��=vyOusYr�l5f� �v=z
l��+���.}�����:��1V�IW.�bt��ş)ϕ�5�&�x�\7V�_�!�?��=tp?�ɏ���� N�(v�S�\��s�8�W�g�X���/���O�?����2�����\,�g韏�������v��s�n��'�/{��ڋ�r�Z㑿�6I��x�q�ӆ��`c��Հ8Fk GDeL%� �N��͜�veWB,4���,�\��`��`Y������J�RtJ]�
�ӐbwL,O^��f�o�TMDSd�^��NW�4iU�u5�g'�[6D$L��>�1ΐ����r	t�3���� 6��ei	��A�5��<����3�`�0� nĘQ�k%[n�8lL����1�<X*ʭ��.1t�7x����>��=�Qj5k=3\�S��R��/�H�8h�ڢyZ��{(xu�b�k�2�̒�P/�/Jf��$���9���ފ��hM����Z5M�����b�Pk��׆��&��4u�C��!֟�o�x*�VVq5Tt�6��D�b�����~];U�C=�\$ݰma���r�;�w/�'L,��T��|����IIA���;��!�9�����[���t�` ���H�޺Mm���|Ǿ��mx*��K�q��Ɛ�S`W�;���6y���M�F
1�r��̥E]V�:�iD:����WD2V�aP�yh��8�����ýyv� 3<n��f'��(�=N�H������ku�A߇j���T:("�r�#�H��V#Ƨ?vn�PeDo�זU�������i�"BZ�o�F	�g*�s��H���c��I|yS<_�`������;� K#[�����S�4�f|�;sj�|7�wi����~��$3���
≝#��A�9�  �Gµ
�z�������D���@\Kcz��7��|�a�9�g�A9�A���w���R�B�)�.>"ؑh�����kЀ��S�&P�uDj�c�x��C��a���^�.hE���1*��oB	W���(q�0|b��i�?OΫ$�P.$�y,s�|t�����?+L*:�=%�*����a��ě�b���!G�Kk�uD��l�A�X� x�ab<^��G�{��ÃF\5����a2벇��Yٯ�][�1����kE���e�&~��JMjZa��m��1�U��L[��b�w���6� 1���p&yA̹�J����^���cI�zg����(�1�S齨�-�������L���ُ0ך�[�Ǭ��B$�S����򶢡M�����AL���v����0��:1����2��������G�{Wa���:t�~�����~;W���7���L�Fv:���;�3�͞��&9���M�g���3����a[}�Em=�HZ�����3�@zgHQ[�c1�X?^g��MS���9��˩��T��YZܤ+��׽�dXD4����%��cG�E�ܱ�͎98�9�+�ݧ�5���s���U��|B�� Ӊs��!�O����D�.k�{?�'�?TW���/�
ޢ��4�̨in�[����q6!T�H+vmA3��-P+�=��t����`��x��s�Y=~L �1��Y%7�{�wxQ�+��U��C:*���.;"�^�W\��RH���CQ~Q3��K��'�%��;�:Pvh�D)#J�����c�!j��|��Yn�k��FE�4��$���Aj�7��Wz�w��9�	�ˏ��U�6���1�K3v�E��]u�mӝ4@R���H�M�g�ůj��yͳ�m�� h����]���p�8��TR��+]3�V���0�!MG