XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��p`��u.���X�e��6�����7��"��C�rH���(�N\eN_�y�ME������b����b#�lz�S�{̓����7��~�)I�X�$������}�*4(\Ԏ7�qZ��˯r���~�#A���Ǟ"�X[jG�!Εxd�>"����	��a(&�>2�30�A�g��G6��:�~Ը�3$�W��d5����E�����A^Ľ1��o��7v�t�]�2t4���g��_�_���CÈ?J鞩�Y<Si���ea��4YkA��(���V�@���ێ���`hN�#q����Be��'��?�a����FN��4���QyY��NGlq�����M"�7��6���,��pb��3H���7��%2P,��0Ӷ58��+������j.�6�w�
�a�?���gN%!V5)@�'4s��sv��ѓ7�M͋X����Y��ܙO����c��g���GW����x�ƂLT{9��a4�C��c�d�H��9�!A ր�P�7�5X���f��ڠ�>��:0�;��0�L(d:��O{���������R�-�#�?ɑ���r��~�^^��-h�?�%����î��%vyշ>7��X�<��q�U��|�r�������>VKo2w���V4�T�Q���0K7��qD�)k��Z�Iwl,ɈSHI�]��[Q��Y��).��Z�`���[B��~2��i!��J�/�ċ$��ǋ�v6ʇ��ڭN��d�z}�\�(��a�6�l�"��N�?W�DXlxVHYEB    fa00    2400�ヘIr�$�Hf��i���0��4�m�\ܨ�a�KTQ頚	zDx�k���я�i�Ͻ,-��A	u@=�7�Ӑ�T���3%"�x���KoE*������c���WX�&P�ݼs�̃Mt�Key�H�>�ft;i�aY.!�����kK����[i����#�]�~��T�� �\yʿ{_|���W*W���T���	?i9���i��G=B�V7�����/<𨲩O_46s��9|fz���eK�5PB4����ӈ�����9������W/���M��^|��H���_Sf�=/AiaKsp�s�	 ��Sϥ��(�������,�S�6��/aV��r�����o����`�LuD
[mI�
fO�F����[|���i��P�����q���'4�:_1�}�UN0H�������|5q������G���m$ʄB���������aCC�4aUp-|
H!��
�9)՗y.M�OpD	���G���iKW�(֧�5��XE9��jJ��N��*�5x��$�4��Ɂ)R����{�X�Y�v籎a��{0�̳Rw�F��~p(���`�b��.\G�O�����`p�0���&��:���j��l���)�HFQ�D!b�K�����
DB��,|&��e�0���jΎk�;ΎbJ����Kẵ���{��	T:Gwk=��E�Rw���g�p�4�Lo�iV�9�$��/�G�!Ғ`#	��TI�r�>�bL��
,�G3�Y�MX5��F��� 1;Q���:�).���b�[�0�Vv�i]�$����YL����kn�LMu����9{��+�e$�X�T?�?�'J�L���9�Q�h�2<���\H>��٧��;��>y�G¸���t���N�P�Vg��[�fj��3�b�w��WK5���;�����N����.9���-��QX)�;.��q��/�<?<%P��6��-7OU�6��gO0�0�/և�x�V����\��4J���������͈���|�J��W%����d(�j�4�Hv�H�AG���+���\ł]eX��.E��������mX�M���1гd�����뽱��էU!�$��JZ�E�0K�8�jA���u�����UU���E.�>�aFɛ�nT�Ӯm�*��)Q�{�i��a�����8_�RW��S
^Tj�A��w*̨J�	�^F�*�/��g�+�	̽W�?�Q���?���!����ޱE}ڮ��Ǿ�U�K�!oS�d�-|�H$���۝h�^���N4)Ii��@b��������8����2����"+8�sI��[rNQ=dm�úM4(��  }+�eŹ��9A���(�)2 ��WA�˟������+�=��O+vr3.U�U{���/�k��{���Ԡ	Cv)!��ȸ�m�5�-~�4�wިPH��<ȓ��9��hS^[̴憰��V5H&2�0�[�U�6�w'8��AXu�7�4��K H�,�֕�>X��=�Yo�Q�<�f�d-+�i��X�v����˩��CI��'Y�}��C�nF�K��f>6..�¾Ӭ#V�2���T�95P� P���)̌���	 �t��|0�k9x�y���^Cr�� �y����Y�u�7|����ʿ�v`#�A?�f�T��֪�,��Δjg��.ܽv>T��`��y ��%��D�ԡ������>3�}y�[�;�N��q���^����Pԋ�|�%',ǜ����V�K,�z�����������CYt�W`�`"+���Вfg�tp��Z��T�A�JiH	�E��_���{� �����Tv��=n�wɤ��g�>�]嗻�rse�u�a��.+d�:6��PjD�W�b��N�n �$������>:՝@]/3��7�����u<T�`�ig\��)k]�jp�+:�(u|a���A��[V�&�:�8KaL���l�5�'?����~Jj������5�Z���Y�����
�/���r&��r�d0��m���Ý�|�ĥRc�No�)�=��@�h��F�/��O�"�9���OB�8�(x�� �5��O��q��:��l,^��7qH�j#��8eQ�2���̑��>M��@3Gޏ�(QT��Z��g*g@b��+��_sl+9���
��/��n��7��0Ewj��ZJAy�䛍d��k�^B�W_�j[�k�MnmY*B�E�,&���x����'�y��+�����(h���N��%���I!c�I+| }�'ʧg���i�lzH��j�~�s� t�������X��6_$఼��p����c��V�^%��d��R��_��j��[��sD�?Q뽥Z�5�ɾj�;BVP�)Uŕs�����eS􏓋(��0/	��N�^�Cn�g#�_$B���~��&�=�$Or �CⲢ�b��-�]����R���q�*b�;p�A�K������v��+�DeW`o[��X�.M�B��>���\բ��=�E�5�0��L�
�PI
�~�
�*�Y�3+�2&6v;��k��M�{tngt��~�l1��Q�G��jg�@'�F�M�j� ��y�|	q����/�:�E9�Y�0�l�'�`}+�N�)ƻ�"i�����Ш�M�$}����/���X�@����1D�-�T�T6�J��H�U��s����S̭�'EJ�h��ů�%P#���n�F�� N�`���
1xu�Գ��Z*Ш�ɢ���� &���x�%����\m� ��:�Ůą����e�ᾊ�&]E�JT�̲[,0og��}�6�ٕ�}lL��}�����Ғ�[��g�����ժ�m	� ���� XW����6��'���ɦ�%MIa�*�$����wi�� ����]7���7�zs�{��g��c=Z�-���������0�'��}�:��f��sT	�π���� �\��`8��p�W��}^�3�sm%+Y�P4S�I`
 p�+t���%L	[ψ��F�Q+Ii\ә�b��;�	ς D�&\u��Ж����H?=���i���C����-u����LG\�$lJX-�}�T��J���w��I�ۺh�Rj��IW��(F͋< �2'b�x��۳X!-��<_T���ɉ�+�b���.�kk��)c���|s�� 5ú*m�����h�P��b>�$^�PKMS'#����٫�/�h%���b����`<H�s�MJG/WK�?�TNJ�o�*����f�Rɳ�$�� ��ޱ���%Sυu�=C����-6T`I�b��Q���<9� {巨���������WkfȑdN�,��������{���I����N�#��'�{��`n
3�>јR Բ�Rl����c�_ ;0�!\���ix�谕+S�L}W
��F�U�)�{X wnr8�M3h��t��&���,�2������?E?����������D�_l�¬s��B���W�
���|>�|<\E�]�a-r��A�7
��+�~��Qg�6tZ�L�d������E�V���ot��l� _ٹH](:}�P]E�	$����;e��r��ﺢ[����V��m���}�O�j�����X|G�tU����۲BO�6��Q�5��,1�$�;[��.S��H�};KY�+5���eY8��Z��b��h�%��q�\��m�����l@�.���:/6j8�-n�p{H��rփ����@�~�%\��+.@��'Ӷ����	L����j����Q�d��(��)�qZ��3�c�_يn/H@׀��#eMn8����]�(+�U_�\���9��hY^�c���S����7^�
i۠��S�ū-�
���_�l�� �̚m��#<���C5T��[�:O���t�
zbO��'G�p��~�ݝ�VF`�>5�s=q_��۷D����p�<�c�d������h�;����N�3���(�db�CG�}���ꚞH�X3B��_�Jt40t�u_�B���;.^�g����>��v-���>^WO�Kd2��ޜ�kQ0�t����g�:v��·�TP��s�n4]j���O6�%�V�t�bٌS<�R\s���݇�D��6�)0r�W���tw�
������4H}ک̔+��t:Ҁ}�4��'2Z=A��<�m2K	���Ƽ��|Hm����2�D�)��7���}	6�M4���;��@n"�{n���P�wǔ�Ad����8�	+�99Let񙁠B�&�j��2�]j��<������'b��1Ҫ2��rS��yDB�0�?"DͬBE��t�C�gbd�ߵhN���SW�00ƅ��H���n�:gJ����n���ρ����tCz�dO��X��@�* �'h����6f@��K�b`�ˇB>~���P���S$��1=]�k�����s/���[���h��;���C����-8�lQ���~���i(T�,�3��M��ׁ� ��w2�:�3p�Z�W�}���$r�Ե��y�M&m�o��&Y��#@d����zt��L����}ރF����JCd�,d�.�ަ[K��{��h/���d�����r��P��bY�U.�P�TSm��<B	Tȥ�\0�[��Ԫ�a�`|���Uw��B��i��"�_ ��	��I�gƌ�y,��EZ�0�9R,�VƋ�Ql.�Yt7�_��'`���b�$����$&O���Eg
����C'q�98���Vs�[� �p��RgwJ� �?����� ^Z���?�:K;��φRz}Zl�&�����{NB\D5�_X�9}��/���q�A�ӕ�T�4�B{����������N�qkT��Rl�(���Z'",�W���U�%[fo�G����;�-�Ŀ���<�ϯ%a�tu=fm�#���q��;�&���2�w�Z�K�X]����_���NS��/��tC5W��pv���}������*\�X�^@ �G�p
�W��F��'�-���P�}S�o�i�w�2�o��om�^�Y��৙Z�I�5-��X��^�@���rӋ�)�Ҷ���D�HC�ӷ]�Od-#[�B:i?!"�O��*�'
v W�	`3�}��uE���M��|���a���ӢZ�}���ϯ��9nS���I�USV	����rE�0N�z��Fj���q�&����|��Ώ*'�՟3�B��I����I9Q�g�T�mu��7�K�k�>?�*�ňm7;�b�.�2� j�QB-�w���=��zT��"q��Y1�A�~&��>iԯ�
�؍	�1���L�ko`�I=x��s����u7ZL+tF�U7�yݍ�<u����?��h^x�;�yET�����T�m6��%��s�y]�ڎ��;��v���v�$��И$;�x{ �B��8E��'��+ƒ$@n;�孵С}vo���z�����[�tc���x6��T��b(��\��+�w4z[TO�N�2�2��>@�c�<đ�x~G��5��w��X�\ ltO��pT	z�d��\/�
w�	�Q�7B8~=d����di^"pq@fG��B��S5b��
�V�mIuk�yd��hn!h,nL,�E�@I���)�=�詌�7�kI�V"� <��VH�gRx�ˌ�u$�2pj�<Z
QQ
WLD��d'�-[��E�ir	6k��aG+���񚱶	h�4a�.v^Q��B"�k��ēmFL�c�Uߖ󡝤�.�a!�(v&Y��)k�]6LZ��ˈ�)�O٬�P#X
���$��X���[x�<��o�Ig-Lˌ�˗��n7+���(�UI;�����0�Z1�/H�
6��F����P�����2L�Z���?���2@>�����.���[Ӡ���Ú�k��$�d��#�xh?"
߈�i��s�l�i���6����^��Y<mc#���:�N�lH�&xd�R��ڣY�Hi2�K���IHap�D�e�����z���c, e��1]�U����I�&OY'.d��������X����)`�`���Zo�q_
�}��>l3���0"{���2��H`?5F8��PZ�-`�B�x��X.�(z�@������B�����0}����|J6[
�f]�[�+�T��~��;����*t9�]�\Y��\�����91j��B�E��hETjы�ϫ�g�ꋃsb��p�7��6I����"S�-�/q[Z�cuo�v.���_+V�?��b�V���'%|	t�8Gp�;d��۔WWD�u5��B)ġOߗ�܆@lJyu��������d7���@U�^X$Tc[���w���*z�a �B�e))��z���"��k�]:�d�+�k/����{���`a^�l��^]id���V��y�'I�DnN�@\���/�厰�l¿;�C�C�/J�m�U,,�f@ޡ%�P8	ɇ�Y��e����[x5p5Koڭ�.��iB7bq>��q6���q.����ê��<��rj<�
s��)�6,]���сD�j�'������m����0�����p����}�@V���OO�>���JdƸ���3=*��@�K�)��C��ɍ:�gK7�ù��S������� }m[�ôR3~`$AF��u����+��PҘ�R��q�-��f��p�S���FbA C�-N�g;"@�1�2�'��w�8n�_*e�p�M��Z��V����>$��/��
��L48�f��J��@�okf&s�O*=<�ن�� �<�ѹ��G%u��t��5�ZU������-.>���}��];#�����?�m��?Pt�,[w)r��ۙ4B�y�˟����p�D�L��S���oºf�#Og0�|<Ejb�|oq���2H� R���}?h�-���.G��5L��Ef�J#/�a�xw�BF��T'���7}��̀��+4y��6˒�d}**�BkTKC/�湎��d��!w6������͊��!�	��S�����Z�[(��f�+B� ���6�d����bgD� v#:9]��]��]��JO=x��wO����Pzɮ�7_��C:M,YB��jZ�a��0�����e�AڟvƟ��n� ck������i���Ք�y��~T��8�*��lØ՞�I�*�o�s�x�8a���򀣳x�x���<s���)�MҔ��.�sW	���~�MQA��/�+j�M��`�v��96�o�/
��Es�<w�J����/z^���˜G�8�6>�S��X����2!ۈ��S��4�ը;�H��m��u�B�� `�g��gQ�G߳G�b����m~�L)C�"P��i9>�@�-k��=:�	^żm44�w��G
�o����V��C�� �;��l9�?���E�aT�i�F�Bx�A��2�%�qR����{�!|���YZ�fUᡲF�~A��;���t��b���b=��̐cQ�k��	���9�[:���c?��ȇB�(�:z�Z��+��^*'=��D�X�m�J���b!F^�^�>������y����(�J�y�����>����8A��ͪ������o|� ��T��xhׇ������x3u��ފ=��C;�;W�¶.u�!��UR�,���Q�U;�=�3���Ii7Yd	:Ǭ�[QJ��r�6�^B��j���E�?)��@����;�P��l�������e)�%�s�{6P�.�����>�U��hN�w�(&g�WVUT��o�J៿Hd$���H��(��3��$+��R��1Ag��<6ma����t��J�)���P[c�%�8%`�#[t��B=DS8��i�%��1���_N%��\���}��-N�EZbVvBq�^��P'��K�O6�.vj��:�d������Q�����+2�JvG�؅-����&w�X�{jnc�;p➮�mdy�Ǭ�:M��#we+�� &��m6}�k���+�H���Z������Ux�o;�w��̹X�0g�a�$�����'��R��u�Y�]�9��JA��������P-�=opc���o{s��o�Ws�ZX�4i��!"�<o��,�bI�����c*��o�)Z��VFt�﹍�rg�e.�I�lS��K�D�<I��۶�V
�"Ė�|�^��. ����L��>L�x��P�6�NX�˟HvZ�J�~0	�T��[jc��K���$.o��o�\#��ءE��ћ���D/�� E�"�c���"�r���3���4r�s�� ���/>�$ٓ�{kk�(����Lۈ{��L\��m�]�{W��aX^�8�	�A���ۭ*v������R�@������=����lI�	�sf�pw�v����N�T��w�=�I)"NZ3%���}��� �?i�M�����^��F�ܩ��X�j�n����!�f嵐n �A"��Xa�w*�se�8�Q�ʌ���M�N�T���#���7��@D�S��t�|������$N��wȺuޕ�R�j��+�5�v���ď���l���C��.�پ�3$�;�<��X���SCd���P��*�F����6�ï�|���p�׺��Z�l�T�ZF��>p��5tm���5q���n����l!hi\�p�x�����!�1)8]�ʀ�F2<����6�t���;Qt:��I)u���8�G��.�У-CƊ��)g��c��������(#Z\�� 5U�:�fr�7����Э���ʶX6��q����F� e�:�^�b��K(�i,�^��.U�s�Վt(E?������	8�Ϭf��w��th��<N�7���긭F�<��i+��p��5_��u�G	���=,�^��i�J�e*k�m�8!�Wb�@��2�ʆ1���~���ׅ�:|� T�[ʋ��Mc9�R ��#y~5�u��av�q��;+n0�X;z��P�"`y��ZX���y��9��q޶2|�XB��H��^�@q���1���gB%���k@���֢GUq_����XM��$�E�:U�p�����������wJ6gD�-㔙ئ2�rA��1�ߎp#У����Ʉ�p�2ܴ/XlxVHYEB    fa00    1ca0�j�F[��ˢ����T�ۧ&i���Rm+&1.���Sm�c�8:n\[��xr� �U�:���<���cECƻ�˳Y��~+�e���޸�L5���F3'[�������g�w�t0D��_Ɩ�� �/����K����h�:� rN�  ��O3F�b³�#��됙��3�b�]A\�[x���z}�h�_x�S'H@� lY�%�e�`�|x�ֺ�J6uq��h	.L�y���t��S�2J�.�� ��%��cAA���6�,�&��2�4�
z�� �c��`���7����'��Tt_�$H�D�m{���%��y�V�`_��Ѧ�6������I���(�����·�H�����Z�Q3�����MP�8S�l�t0���*DY;x�l��ڣcˎ5aB.�n��4*�;N�n��F)�yW����l�}��}�c�3����"x������>-�H�G&ѭm�'J��VT�T7�memh�����~����|�9.�A0,���Gm�֌Z�5���R���z�a�����Wl'�--��gx�N����� 5�X0�ԇ����A�t牕](�`!��x��H���d��:izy�b�v�7`�.�,[.I�R�㱐  �#�{�}��%-�n�m�t·��=oܒ��Է�(�`M�#o�v~1B�Z2��t ���D����Fu��^g/�P�N��o�U㭰eaĄ[��3J�Ti/x�=ڞ�5�3�BS��D4���K;�8��A��n��O��`~Й�(A7�6'���bH�[�2K����3�a�M�S$�q�f�r�?�[Ƅ��1sP�-���L�Q�<c[6�`�.��bN�1p���,~}_�B8��>+A\?��1@B��c�bv|%��]s��`b�ߚsw�r�8u�fËJ�RE�%�g>�
=p���]�j�OQ�3Ӓ\��!�$`�2�4��F���E'�Z�<f�~aB�af�,���)Տ �;e��1���_�	��漃d	��Y�¢vቬ�ș���	�e�4%�����mo�BT[�H�ޣ����oA�������
#�U�c�kKCy62��I�4d	�jɋ�v	 .!]�YUbt`�n�ɣ�!ќ4e��5kl�߳t,Pk�{�rA�)�,�`��_=�5iA�s0�m�V���97�c���|Y����Ȣ�	I������V�;�Z-]{��kL���e��
��*�C�n��lՓ/�1���(�P<I5�eڌ��	�iӸ�XoCNSE�w�"�Ya)%��|��;R龪!o-W����i�/��u�
\��Xx������. �K��ͨ J�{�Nak�>���S���J]a,��!s�*L���cs�B-WMth*���m��w����������r��6�3�����}��I�@�[�}�QG1���:u���|O�����5�b�7� ,-�`0���>2"�����Lɍ�s��Ѹ����3>p��6gz[;"3��&93>s� �ZV���,En�swA|�\�N�*���+O.��g���H�W�3��U?sS~�J{���k��#v����e�\D����E����LՕ2Wy�5C������6�c͈X3�Ȓ'�%h�\�t��u�F�*U(����ܠE)�K�O �kԀ��+�]���,�`m��1�C�0$�S�SW�-��x�_e��d���t�!y�ˇ��A� S`x�*���d��r��F�������d�g�t��ഌ��-�!A�����C
mgm�'��k[��Rq�7�F��{�e��V#�
#n;��V�j=</��N�D�.T4n�9�N��3��N�h@� �z�<�f\.P_P���2o%Е����P�f� k["~�u��;9��(��k뤝!G�p��d��k�gB��_n�7<����K[���xN%�ۀ�N��H�r�\��+0GS�t�slw�h�flۼ^˅�G���L}X��[5�\�}3\��(E�>'f���_�t�$���.ڡ|�57�Sr�'��,��ךAQ����#	 �	nd����%;L�� u.�qġ���}6�x��Ž�h
C��UY�+�`M�)M�����@��.�e���=��?͝�))�:�@d��c�`�R��C��]\Tp񧤆�?�;�~����`]"�V�"���x���;��{��Y!�>(5�щ���m�l��N�ȿ�BU'��5.B�~�࿑���
�m�
��xܕ%�� ����4:�9�bS� � ��L-CF���A������'�2���H:��,��r����G��ID���~��=H������oI%��a���"w2��9�:������4u��"�׈����P��ȑ�I}:��7Ia��䝃��U*\�\J�b�zޖ9j�D�Z�#���4�����BOxZG�$I��㓻��
��A zI��q�R��PփvF#D�bZG����H �n/���(Ny�﭅y��^D@"aP;DY%�oyd?��U���OH�i�U?�<�Ν��=��z�3v�j��$%�8�.�f�����=���T��ә�Q6��l�)d�Ͳ�S�@��k����y�@�_�Sϧ�r�Ҵ���y_`�I�%�-m�ҪDQ�Ȱh�0A:��_��#�4K�彨�GK����:&=m�"9~�*H_�[X���j���e9����i����L���I�����裬`�>V&�n.�͎�\U�	�Q�w�	-]��]�u��1�m�%�x�.fYl#�Bl��U��j��p	�t}��lق��&$�0�����骖���<�B�{����@����Q]����T���N��ߔ���i�+1�#S_��I�Qe��63� �u��!u݅�_�_���
�\,*3���L��㭹T�өd�J �r.����N�[ڔ���/ �]r�Iޏ��OY�|��ȭ�	*�N%��R��wA�Shg��sٔ���sR�G�'�&�8�p�ݶN(�\Z�t��8�p��n���ckq	����i�4?����"#�6.�����.х�'���?7{��)K
s!_&F��%�G>ّ8c�ѕ|����[L��3��H	�ѩ�Y"�%���;�D��Um:�}��\���0`,K1�D���ɪH��E�{u�C��q���Ӄ�N�;pl �����t^����zt��F�	������F��n�6���bmf�{ge���6JG����^��1f�G�~�D=_�\5�[3͊K���e��Oڕ"/�6qo7j�5��ݏI�����KC����R���Go+==��0�{v���x���x_�t2�dX�E3,<�z��"�	�
�)�'��h3K�-Ϧ��~�<�3��,V�je��7�	�J6�e חi�ݎR�ڹ�|����ʃK"�Bp\�[ʑ޷�A���p�M59�޵���2V�՗�ŏ�Q�.mC��]��F+�3p�D���q�d�J�����>������9j��#|�Ƨ��@��-��At",�:|�H�=f�O.�:X�~���v{��l�T�k�r��ƭ�b���T���|��|���ʂop3�_�*�����P�t�5Y�����9�n-�'b���z�;�4*hp�	����Q�`����w��nԳe�4%��6RY+Q�龍=x��\�x����ɐƇ�ʆ3�_�p���1eaA0�g��MiW89ߺ:�4t����v������	~�&�s�d�����V^���3��f�b��C2���'��j�%�zO峏}��ެ�= Z��+^����,��nB67�M�S/*�͈��\B*�c����ښ�~3��zS��!Y\�C�E7��LT��:��Q�b��Du=���������1��NBMv��6=Ô62&���{5MA9-���ï?
�P͓_��Y�4���.�DӾ2:7�
N�|-�IQ�\t��\�S[�;r�-��v�A��\�RE'rz7,2��%a����veNaff ������	�O{N�8ct�՘h���$�<�'�/��c�/+��.�؇E�����
{�2NSC�D�U�K�����Y�&f�(Ԫ_k*��m�v�;�-_�U�8�%:aR��)��B$$&�F������M��F��7��A����`u�a�����A�i��nf�˽��W��d��yr]�ML?��v�Y�\i�Z,��^���,0w��$��� ��lxb�tN~Plo<S<���:�э�~-�	��7�p�+A��_�
wp
w͟2R��Zh7�=͓A���%�P�{I��sU�2��P�N�ZE�����Y��{9+Za�;!�gq�tBA���U1���M�MW�1�ud�'fAh�plc}��5n������*0�-!��2�������2��"���KY"�>$�`�l�>H��u�:9���|p/����v��W>�k1kA��S{ u��_B�í��z��_��W�����ѥ�����j��5��^_��+�C�b
�>����j��#.f�ɭWy_3;M~��l��G�����u2��ŷ.^���E\�a���ư�A�^3�����	μk�#�%���AL����E?�ޣ�q6��5sǗ�\�x�13v)�i����OV�h�pʮށ?�/�}_��	�;nj�1�ܰOi�=Q��a��?�¬�;��6�H��Q_s��º����E���j��8-v��r�����?�ܠb�7>!������i�#�&��r5B�e�[˽K ������&���S�hM��ܻEP.ɋ�w�bk��'��>-����>z!Y��B�'�>�'fU)�x�`A��Y�����������Xꇤ��I��uM�<xE�4���_d�O<mʜGp��s4���[9EB0���ŊG�t;t���ߪ�>���^b9�_����
����ֲ$f:��Q���=`(�`宖���5഻��>-"֖�:�]k��M�exs"�E���R�deN�jf�.�(��HGB��:�~ƙ(�P��S���I���#:I�m���|�u�!L%�1��ٌX\��u~6������KЌR��u�*�~A�@��:��d���-�'M��B�$��Pe��*�-��x���{��i�$�z>�%���=>�뷍ʍ������#��r��jU��3Q�m\E�/\:	������s�#�&�Q8��t!컂���Rc�D�ǣ�����^��pÎu�k4�"�!�#��lMǚ�yϖ�\n�{�M]
�ؗf�����X�a?~G��G ���n��1m�l잭���B(�����X��޼
M�������m�ۋyW2=ۚ����ݕf2�	���2p��k5��2�q�,��4""pV�p���ۿo��6A}��:#�U��T��������ۇ�<!��+�������9��m�(TU|4ϕ`�:̆ٚ͘/�T-�:}U��<��"�!Ė�~qϢ���ʛ�rz�[��&��� �n��S�w	Br��,��j����G:Rk���)���P�\�a�?.�ee{ϖ)3�e�$�/�~��
z�`Zǘ*򼓒.3ԡ~�)(�/�Hy��'���膏{F`������SAY��=�K�qNd��l<`�P��}�}L��%'�YHATj��wE�1�7{	���9�K�ƭ4�OJi/�G�S<��:�r�f�e4i�Sݦ��BO��g])ޒqyԬU�O��s�+	���?�n��
�B����ܪ���=n��#
�˱�?䃂�q0�8�$��7�h��#@�ME/�p�0f�pK^×0<oӱb���Ϣ��i��p�(b�N�p��� "���?��'�����?OX� ���? �br������5�&�4v����m���]T�x��K�CY��H����^O>���8s\�����Pl��[���^����^ob����Q�(`��-�-;�.ĕ���p��rn&�"��
�O(�.V՗=Cj��ǹB�sS�xo��F�}$;�i�2BD?�}`TtD[R�e:bbG��E+�F��?�'�,�U�����L��<Xq��G����T
�6�g?�u�|�3}^~��48���K���AFE"g�k/��SM,4w�P �2�J;\b�s?�nϑۖ{�s)g?�嬢"u�3����u�����̫�G�WB,���?�gm/J�[z���7� ��=�?d5�g��=��T���.s�'�Q3���]��
+�W�+ܓbt��=�X�A���Uc0�F�Fy���K��\�4�cn�?,Q�Gw�N
�k�(��]��Q�����}��v��D4*���1F���]�DP�\�@&f�T�Q� O��N����V���}�?�*���&��T6n�q�-������� �g����d�Fe���a㛣T<�g�s�n'�_��
s�/��)_��ŭj�Ûb���(]�nC��@D؟��ߍ�|�r�cka��91���\����Ӂ,M�����s�Z*�Z��'�m��c�A�i�0k�Q<��4��|�R����I���a=������4gt=���y�7)������+�ܾ%���`V�OI<���0��*F
 Y:�~�{)�w�76��aRMOy�O���;�x�*�n^�㻚���`r�k���I�rv.���hۍ��'v ��W��߀0MfE~Z�v~�^��?��"����g.1<�{(:G��G6_@�,'E$'�
L���?��@�H�X4U1��&t5Wr���tZ���6a�+�p�3�*:�b�F���p�s':~�j��s��{0�ͧ2�g2����<��t�w��;����ထ��1�Y>4�
��O��'��ǎ`�~X�D�v[��Ԕ�sE��"N�)oa�څ0_�Wpǉ��/�1�Vp`�Q���?�~����m7`�-&�u�$/H�����}�QR��<w�NWL
���km{f	�[&k��/�fS�O;mY#*z�:��MZ���A2�m��f�8Hd�'�&��1>B�R,P �m�a ��{��O��?�&~�ĎVL)�V�?�$�q�P�"93���W 7�Ύ�6~�v�q����vac���g�F&˦�0��@WW�h�`�8�64�s��ؤh
�<t�*�{�3lӵU��<�.�bXlxVHYEB    6b84    1270[�k �oY�{�ɈU7�,�L�E�Q_�E8�\Y���	� �d ۧ>$o"+��--��//}m: ?�}������v��&:���3|�g�'F�[������(�>?Lk�*}���~�;��<G�q(���ݍPK�єB��k(�^:�9�<	e��L��S#���4s<,�q��e��T���+�������0��x��������vB�x�<Y=�U�}���~2,��>����� �{wٕ@9�L^�c�	�4nˣ#�����|Qr�W�xw�+<� �q�b\��=�B�^yI�f�G*�n�D� �d����D:W�<�p�^H�G�]�M�����Qs��n��|\��?�Xd�K����f��	C�<E�� ���l2:t�KQ��M�^���IʢQh�̓[&�(�I|�FF0�-��@m�V~� 5�ZJ��V�m� a+��ui���F(�	e{Bc섯'Ѭ�*%�L�kb��-.kle\z��RM�:cyO���І1B��/�i��r	���CBH��L�iZ�:��ߐ62�w�A�mP	�)��fY4!�-)|��O��d�h?�}k�Vo��#���zG'�+%�:$o.�q�0�H��������b�0��I�2���c.P��ȹH/{K�����Z�O]�*�]?�ªXHQ�=�xu��_��.���#1�8q�� I3��tË�dW�ͪ��G�U����m�_gBJ1��� !����{+t6��$�O��ưo�p�I��-��Z{��MV�&1}����z{���M��E_p�yL-�`����.(aS��3��k~�p�<�R8Lv��)O n�pQ ��C���BԼ���ˍ�P/�� r��:�Y#S� ��" ^iWV-ꗺ�x���K�2�q�"����{G8�=��D|N����\& �B�u2v��)7���L:�@����+AX�0����t� |�Rg���Ι����D��ػ\�0n<8�\Qv�Vv��B��п�Q����	�N�6��x^{HZ���.�}=��V�����Q	��8
r��~�Hː��'vS�n"Ɛ�ţӍ�6��Z�I�Z�?�9r�:Ҡ�mt��p�"�������䯲$�BJQ�!^X��lLg)׌����P+"����vt�^�����*$�8r�L� � ��L� P�M����=^vE�d�>��*v�E�g%06[�>|��Y�H���;?�'���F�}����s��"��X��'�,d2��D ��4zA�_����f�2l��Z<s���vʓ�Kߵ�d�
pV��N���~��~�wg̖k>-�l�F�{�h�W�՛���.��г��k'�{���9�W\Y�|@1(�ƽ������"o.�aJB�6f�J���c�0�7|V�;g��KJ�Oa���l�~�YCf��!�3���kV�5)����$k;]�������F�h��7�������]�h� ���]�F���΍��"�3�&��K�̕B���Q8E��D�����9L�����~H�P��2@�:��-���gOx���P���&m�d]���o�$ޔ4�G�����>��o6>0�]�[M��(�Н�}����.��u�D{��� %��ז0�"���uz
�Ryb>ɼH����s�@At��Kn(h���l��1􍖱h��������e����90�g��|Z}����*�q�u�ʬ^��D=��S5��j20�f�4[�t�A�����X��6��p�9��y."�60jt�VP��@������klu1u����ޫWF���5#5��t|ch9��W@�~	��j��e�osG���N)kY��+�Y^#Hy��P~�?��'nPDݿ=Gf>�6�X�Y!��F��~lZ~��������>c6Z���v��*�9k�q��H��|P�QVKk��o�vvv�xd���MD�PE}k�q<%����㹎Z�_�r�o��7 M�WEf#/�9�$r*<f􈸓�k��xV�_�X�f� �ol�RD����&W��Җ�EV�¿I嗋�wJ[�R� N�6���+j�������C5����,���K�}����S�8>���̩�?d���uA��}m�\��)&)2�gB�����`%�p�|P����|�q�!��%�_&p�I�dg��(p�����T�I��Y���Xo6�<ե�o32��C�We���Ƈ_�����G��g��Ë���wz�6ʈ6�lN���UJC�p���p�2�L�Z�_7đ���8�MJǀ씞Z�C�술����Iy�^1
�V]�K��{!����);����_{�9��[!*ȥ0�>|S�*c�����������z{�\����� �@Tާ@��x��Phs��jv���i��k��ҭ��*ا��v��$]���pH���maL�S0^ؐHb�?Np����*�xh��j�x��9G�Yf����5��ʘ4u0����(�gez3к[ddB�n�#��=zG.�Lf=0ʿ&��
�ǧ�l.�y���������a�z������-���4��������J΢����vU��t�x�43N� �0����×����������I����0�����5H���/���:��|
p�{$�H�F�y"��3��& �Osr»%�t�x��>�~�}Q��l��_B�>X���ʯt�(��D����1d��m!�س&��˹Liq��m��%!��tW*�ǯCP��c��4��x�	�5$S0�۵��#�;�Џ�0�E���-y~�E��{7Y����D�JƑ���8��O*�A%�ׯ�G�a�4��ځ�}U)`_~(����[|}I���;z?��\2i��p��ܥ+�[:�r�YJ�q����[ϔz��O��a<�T���[�P8�>�}�B	'a�NE�t���`<���7ι#|#�s��m�&,�R���C��'(�ٹ/e����2?�g���G�\{��$��~uOp��m��VHR!�oe��ܳ胠
g]�FU�ΖT��_�m;t�F�yjc�u��Ƹ���\$v�|�y%/��H�=��Ԇ�]W�{.[�C�N}�`�<��ߤ�Ɔ�q�7��y=@��ùhm��G\T�t�92�Jl���,e���șNBob�K';�'��m�6��Y)8�Nv	ධ0Z����'Ph�s �64֕�ެh�C���sY���_�~�^�;����zS7����o3�!1���5*U��p�zg[�j�*����bUٵ΃'w��<|�߻�|?D<�$0����Jm����AJ�Jl���7ak6?��U�#�zR�"��Pq�{&��SL��,"ݣ�[u����,����Z>\���r��rK�z.T��s�1p�J|�oW�*Hn[�!x@���V�·���Ӱs�HךG�~�E%]RZ�&�A�A��44��вCR�̐xC�)<D[_p����uE\&�������L�Gp�	v+��?��g�M����gfi�J��
-�/;Q��%f>�0����0�v~�.(��:Gk���O���*���:�D��d���ыGzkL1C��ָ�OE"\i��S@�DHd��EUn����sZ�!�B�O�0����G�@�8�1MSX�d�mR�0'+i����1�ȉQ����n�b�i𻧰�s-°}
@=*�^yX.~z���a�+)-��L�;���p���S�����\f�<����
y�_zli_*��GF\�2+4��y�Ô����#Y���E�)��8��
2�f�2���	���<���5y���]��v�s�!�&&H/0�v/Fק}�ܑ����i*�]�!s��/@q�A�$v?V�j�;�u�e���N���x�q�/�gu���{j�y""������.)�V9���J�測NW���4P�^�&_�%�ZP��a���V��%���%����{c�p��۟\C���������#��Ƨ���.eq;����T���~{̷�
�*,�sb������xy�����}$FX�L����/l�H0��� Ƞ^�hpT@�.+���<ؗPj������X��e�?ea�-ƸT^'�żs�����3�q�B;� �RZ�I��[���B�Ws3�}Ũ�<��m1T1D]y��h't�G�#�Ι��1�F�>����zˋ"�ڷ�+k4� fx��~k��lU��I~khW��"�U�q�w,�0��*��6`G��S�r@�N�HM���[�����\�x�R4Y�h �2Q/��W���Z	o<*ì��\�{7��i^���_Z֏Nt�3t���l����;�(�\������b�,���ۗ�ˣh�(�t܁ĩ3���f�J�(���l{)�APWs�e�� ��#�W�d��sJ޿�:*@Q�k��,�TtIZ�����pt�l�'T$�/����Ϋ*�������FD؄��
+|ӛx|��j]s��̅>C~���;C].���omb�1{��	?�__D��p��Nz!����de����j�?����}$nsX��IH�*~v�Yݘ���Ds7������+�{�JY7_)��셃��@�
�@K�}K%��z�*�o��U"��W���ͪd:�xe*��Mo�b�g��8u(hmSm�����=��W�