XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Ϛ`-_6�D���ח�`ID��x)-����]d��M`$�ʎ@��@1r��-��^���
,e�
*n���<k�D���Sq2D�?AI�K|�(%x'ٗ�@ O��Qo5�0qX�-!#DIWM_y1#�|��&4I�p~m���Y����n�G��j���u�����%��[�`^p��^�Jr:��/S,]˙}��?�q0I�![��̃�HKq�յ���:��Dh_�=��������jʮ缿�B\�5�1ZE��s����ӕMՑ	������I�^Ce(���VcLd8y�p��@���Ϥ��]�e��( M�BSAgұ�2ǟ�n���U�G �>",�XW~�h�Yک��&�����.�|6�� �2X�7�J%ڟ�B�S�)���ʃ.���i��_�L��Tƹ�ZM߇q&�����q�� �a�lݒn%�G��t���0l�hm'����L(��N�k��^� ��74H��������m��'L��ݾa�T�z3;�Vy�j[���%Ȯ�䰆�����Rw�B�PD5�S+�z[o�H6��k=C�8�v��J�i�Ns��z$�'��������WJgW��v��ƨ��u2��B�o�w����������H������3F�v��j{'.sS��ji��Erյ]f����p۝�Yݣ	%����> ��o9Yz7�
�.��M����?�.F�[Az���@j`�`��س�;L��DɆ�9>�=D׌��"���XlxVHYEB    fa00    28c0n�^ږK�"i]O�/��CP//�q�R:#�U8�Y���E�k�%�i��pU�����&�x'�w���|Xu�ۅ�H��(�W���z�Q�:<Z@����QaL�C�d4
�7���U0��C-�`ul[u`�����9eWۈ���]\�7yk��c�����,�R>��H�,B Nw�ؖ5��I�1��iZ?Ou��`I�����}��y������YrE�zFGie�y�.�YP���?݇z��?�>G�;�ı�=��A�������h�j�^h�Js���,��|�6"�\���p��ɧ���f�φ�,���Zr�>�P�2j����\���a�M@�h_!�aO��Z�KR�Vn(�(A�T0< ��be�M�93��!
C�͇VNDC@�"������6<��l�<�T�p^����Dx�<3�P����u�ǲ�PTɬ��f���[���g���u���*?Y�2%��	��&0ν��q!�mo-cʎ�e0(�1ټ��[HLJ#�r:��e��&<��ֿb�V����:ʴ(t|�
p�W��

�j�r˩���>�v�=BjLQ�U��=���ߚN�"��g/:��"�*!v&�$��VE��0TL��@n�i��H?����%��w����D�����=�E�"�"��Bʆka2(�H�%~^�^�����JJwث�$��i�=>�B|���@L�ڃ$ �up��5W���������r���m ��ÑX��@Zc�N�M$����ΌS�.��p4�9D3��Ys�l`��r���>�8Pld���3�%l4�|x�7G���$�dP�vr=�bF�Z.�K�+\un?$���OD��а��]ZAj.q6���7�ʟ{u�e��97�^5�J����VS3�K���*���9�֜征P���t���,�堻L�x��cs`�1�8�'�N��1<��=�1�/��!?��e�\+�y�����)�F<�׶�����(��S[�,U��Mj�����+!�?JN�CEg�A	�)�,/ )�R�6%_L	��}N���fT��>
A�r������f�ͦ��M�,JV���E��s�5��SԿ�8E�W�W���JӞӏQ��GGD��PѿpJ�h��D>ɪ�2Rrt���45w��}�~�QD0��ɰ�W��T��t|@��(�`1ԛ�<�R�*S��ѫLj`T.�M��IY?"�$\%]V�GL��UH�]��.��7B��B�8�4���4����g���t)���׌K���ܽ����N�u�3��2.8|܈��]E�J%s��쫖���·��BK��������-�y\7����WB�	 _�>&���d���:1�����!~ܩ�
�.�GM��)�BY�l���A�B}�_t>�tT���`sY%�dJ
)�x��KҸ���r��x93
97*C����ٮ8.�hH�Y6��|&�R���c_������A/z�':��679���M3X
 �0���B_pg�=Ʒ!���h���Uc)���V8#"�diB}Ȭh�@
����8���S��O��7�����;UWg�Et�^R7e%C��$��@Y"�bJ䤃���Ft�DN��l�K�����'+�4$�=RU���2��x,E��$Y���A�j9F��ʞ3<�^���:��ЗR� %�KP�T>�����2�d�ԳS�1'q�T���8�k�H �p�P�����17͐�|�Y��ڤ�{$c�4l���5UTj%��I�k�yi���U�oz�-�Z\?�Z�Ѭ�����s=j]����=K���>hX�s��j�g�-�z7_�Z��
�)��SG�m���g'����PĂ���)�M�P�ޡs��M��C.)ɝ����Sl��ף(��P��-��I�h��Ք��|�%��ӑ]�<�YU��u��V��IZD�o�㨿@AbE%���Z����YL�^ d���$K���V�=_}hP�rw�2�5#�#>�k�'�^�g�/K�������e�����f�JD�)^^�i���a^�1K�[@��������>_���J��>P�=�_)�$c�䆾wO?�P��f��C!�Y�dRO�P�Vk�&��)�h���6��j���SQ�M�}� ��p�j������D�z+��S���Y�$~�\�5�θ>�S�'P���Z������M�=[��8r?H{|��,�w��""���mHe�*18�"+�O�_�}�.<�J����W��'e���Us�G,&@T�%`��$�ܕ\ n�^���\���C���*]�W_���S��_|���Q���7%�a�xR�.T��̡�C���LaH��������Q��.��	*���D+9߯m��T�lV*��^!���;r�%�ⵈ(�8�g�M�L�p�,G�_��f���jR�w�\��D��U��5����k���|�㧦i�3:}L�?�S_U��Ǘ&wQ��PR?��tQ/�`�9Tc��ݖy{-�
�6*�_�L#P��j
�����B:A��R���Gj��NzÐ����·C	�c����Y���
`�e�/����'h���K?�ꐢЇ��y�����n�y�U#�[���Y9s5�)�E�6C� �)��8�+�,�����䕄T��ՀzK��]��}�Z��a���C�&r:q�j���Q��iQ��p �Hl�P�'��o���u���s��i�ݖ��Q�v^�p�(�Q��	�����kA_'�[K��׊��p<����f�z�w��qXg»���E�O���^ҟ���CS1%u�u}��sf�H��n��d�PjtOZ��-C�q"kڬ*�=����E���'�h��q�}�Ɋ�(˻e�n���=Tj:�3>�$��
�j!��6�8�@��B��q� �"gx�j�%@�e�pI`w5�)����/=~�ϒ��p[�C4�ʞ��kߴ6sn��+���ej3óYJ����"��G�v
#fL(�/{x�OFfZhj�<��H��׷��b����1�2^%���b�K���Ԧ���AL��h�^�`�OC�\+ۈ-~�N/���$��tJ>���Y����>d���eq��a��b�F>�K���Qn&v�E�kŊ����a�=���1��ڈʇ[o�ǭ�9�|L��w[��u��w�%��|�?���!���kh�A�~Hw�mH)!4&��k ��l1��$���&<K�y%��8,�1͜QR��¯�p}��D\1�U��wZE�i�V�{��0��\��5E}�����x�Y��)��*���y�S���B넹_�@��^��#��Y/4�4�@c���/�����߀,[d���R�)sf+)k��o��"֑B��Q���n)�W�uʇ!���s�j��h�q�p�L�MK�������]~�x��`�-@@5���UM�f8��#?��2j9c�ym��d ^V�U�b��6)WR��*eL8����w��ir����Z ,��b��+�^�xP T[��.F"����W]<Z�y�����7~�(Bq�\�X*���B�h&kRZ����3s�uB����	�ջ+�h�>Tj��!�D^�p�@�T�=L����a(����Q}y�߂Mt��U4mK���(�b�+�E2&�?�8�Y�0��M�胔��b������xh����X8n�T�~̱+>�%������p=b:������1����ԓ���v~�b��"����徼�n�.%�+����d.�M���@��tsծ!t7T���'[����!Yx#�r��2�K�`�El���������3����i	*��Q�G���t/
8r,	�2L �M�U�k\E�N�����=ΈF�T�fkug�q�$3��^r�v�z��c�mQT�%��͐�qO�����`ަY��� ;�β�imqB�2�L�����j4M߭i��R����J#`ԣ^P�����l[y�/-�l�Zv��2�\���8ю��OY>{m��V�zHwv��:Qb� p��]ڈ��u3 
=��v��Ҏa.ڐ�g�><�V��$�(���Ե5��Ԛ����O5� �-.Y,(�
ޘ�90W��y��C%$��C�����g�E�,6(�@�i'���6o�Sյ����������ݍ� ?S�n�C����P������
fG���A܌�+�Ѣ��6?��~�ͩ�:��)����������rL��s�nsہ�
7��_h�|�~,�����7^]��9%&3TI:��/�H+����,7�/� ���Y��&��2�~z,�����sW��"��9���F��XX�^��&��d�VQ*�5�EAc��T���մ6���G�é�̆Z�V���E� kXN�'ͫ���o?�h���>��c4m�[��<���LԲs_[���|y���_��ʪ	Q(Ot����˲<�<(nP?�f���J�_�^�/���7xu���VQ��Awqm%���ސ鼪]|OKl[3��f��!���y�&R�%�-A��ipH�sӊ=�Ru����g��3��=��{�r����a	'��7/݉-fx�V��t���(��w6,= [�������"�3K�ps��7�`�;Rl-���r��v��_s0�퇳�1'�8�#�6��@�d)��8;���\�E�	�MnE��oa ��OBĖ9��Z�;�C���,Lt�M��:w����w�|�:�I�C�7�O��@�����vdvGJ#{tjG<�o��{
�L�n�C����T>����	8�]�z^�x(�
�g�g�2-�����������b'RP���h������8؟Ԓ����H�Ƥ�s�hF*-�a���-C,IŦԼ��U�fi�;��V���*7d���U�ٞ��R�q��a��w(���~U۳��-��u�3�*�,t�Z��q9�Y�ѫ��-{��yW@�.?;�����y���ysr}�fԛ���j�:k�>nv�'ni����]��D�!�d5P��wo����|����[�;�n�w����#̮կ���M��u��iIg�=�#(Ҳ�Lf�D"Y@o}*��K�= M��bc`�v>3q��=Ԃ�C�t�;�ѼSgS��7���p0 �?���|-ZK �;���n|���eZ;E7c���=p�R�)q�mU����.g��6�,Q=����ὣ]�,�F\�Đϫ�ڋ\`F���n"���2���L-�X�E�yVy�bW
�^��z��#�a����"n= G������V2������$D���ڒ��]�C��=���|?�=���8"4���Q"���V{��a^i_Gu��둤�)�$�h���{z`:�O\�d�����g.�J����|_��\�9�Դ��އ�5&Y%��K�o�QT�n@�/7��;���Ϳ���A���Uk�����)�x��Vb�[���&T}�@�n��D�*$�X�WBj��?��p�S��9�~��q㶁��(U0�!���%��w�nq;w��U���a��R/���7Z2�xBv��9lB.�u�M��^&�/�~��Q��Q���斑�BEH��ʡ>��v�W��EQ_��UĒ> ����}��
U/�E"��$Ƒz�ι3�l�V�#�$����{�p��J%>�i	fXCʚ�d�Ќ��3���C=��A!Qv'�� z�`ꐮ�	�Q;����ㆡÙ�)5���>,U���t�"9_�q��	�h�q(����M��>u`ڞ~DYDx���ԅ	��2�@�#�1P'b{�iJ�L9�R��?��Og���o���j�'���I�w��� �����$�_���e�(��H�I�+.�]�7�.��b��h#��a�`x<G�}��w�������rT ����`bVI~H�c�w!%o��^K��3j��ꛣQ �{벌�,�P[l��Dk��w�S�� 6Kj�����&?E$ɉ�m�t��P�jj��.������|�ٸ'п��nь9�UL�ہ.�T9v�TZԑ_�6�����lh��ј��71�|���1�+LndI7���I�K"�e�OY����<0���q��S�h�mO|��i.
_W��~���*�$j
�́���/R&Ad���WC��r�*3Tm��H�3��@ɴ�j�"Cc�fgk�6;0cX�z���*e�K��W���u��J03J3_��OQ��tn���l��h�*������)����߱>7\��B 8�����p]P��ë?B%��}4<y���L�~X��� W? h���Wa�(�@!�vJ>��o_t�C��H%Z�=X<#��S���4N`� �P�H�����J 1����P57�?@.�;��j+�
m%�f�]�W@{,
��ߜ}ُ5��^X:���o���KY1�pl�ͥ��.[A�oab��fx����ƴM��:�Jl�S;V�}�c�$�����%�����J�`M�粧T�e-�Xã�X�u�m�)��_�&1o�g�t�|��}%>�Ҁ�$+A��{�e㯓@Tɍ/@#�b�{�J��Z3�8�*�V�^Bl�&���g�>�+P�_}��pj�q���f�˲��Bhl&���C���e�D�2�>�i;���:�!�pu(�]BH���H�jo���/6��
�M���B�
��m�d�p��$����QX��8"��18��u9�}���o�p��x��eH����5��XT���3j2.����g1���t�3��q�5ˑ��;4TB,�{���0�S'�K���hU�<�~H|-������WUyƠ��as U^r��(��<��S	��+�����I^�ֳ�ev����46��� 4��nPg��.��>��K룷��q�c}���u���s^5T&��W^���-�L��!���?y�p��4a�b��ǚ>��a�ʋ�5j5ˆ��P�$^���]W�
,�����m�2����~�S�\LN���g$�}�0l��7⪹)H���S-�w ��W�3(}���<'.�DO��9>��9g�#��w*q�f���/8�ʀ�������s��"О��^2�ѵsF\jsO�K �5������<إ�\_�~`�CD*�-�2)�Ӻ�}��9t U]�3&\-#���}����p��w�����H.񎆲A���e~T�����֓�7�#�w��\|�I�ܢ;�!��aXL�a�G�%�ެ��A�������g���j�!��������K��O�ֆ���Qp�p��J�:��y���ސ���ٍD\	'�%�_y�?Դh�WQ�jxè
�B�X��URs$e�	w ��`\H� &H��:��䌅�H�e�.T���̓���aZ�ޚ�*�|�z��R��m���<B�H����o3v�lIi��x��#�tF�F�u�����4�ɉ?�I��?��L�(N��o@�@+��w�i�?� wI��$��6.Bȧx�m����s�KNƀ�Ջ*�bRK�����r�`Fl�R�vQ���>�;t��W{��jp�^�3$["��vx��J�4��w&uA �mTH\���H42�9�B�3�km�T�S7n[�{��^FM+F-z���s��'\7Ήn�lU��'��I��~�2��o�qO��b4���M����)�Ql�i�W�Ht�l��������unÚ��_@�ɓD���7��>��,���h��N�Y��z �B��'Y'Z�n<n�!�']�,�3w1b��9D�@�^ަ4�4�jUՑN�>ڃ�p�n��^%3�QT!P�m�{z�'\���,f�BWת��{�j�;��,r3�dɉ<�!�ߦ�96���ض7� �ڭ¤Z0$�����Y�>j��:0��G�t�������Tt1!y_���akR<zҽ��,[/.��Ġ�� ��!�)#W�\��;j�����8����ZG�wo��WPݴ�������Q5�
�ۯ�`��IɌ9���Tm�>��f�3��-$~�a�3,Sq@*SH��\<�3��q=.�90�f�x��C��!6lzܿ�����h	A6�N.z�Q|;?��%�b��e  �UB41r�`V4��wF�%K�O^�qX%�x�{�ֈ9<T��y2����Xu��gޱ::-�{l(CF�g���������XiV�e� &�s<�O_�S��k�_�u9tV�����5��!/{�bБ���ş�S7����9e�T�χ�J��(11|��Д�J5�^jpz��1RYA=\��}��G�� R;d6��:���F�c�jo�EȲ��	�>�������m:%E2 *$�w���S���DV�¥[�⯴1���i@�������z\fD�/m��q�3[6{WH1݀�-�;��X��zak�[2�L�]��u�Ia������3W::�ہ��qz�Ep�M�RCȳjJ�k�C�~����*bV4�(�@q;2g���������3d��	��k'�&fC�W���T�F����ч�_�-��r*�G���o.fJ�xgXL,�!]�
�LE�������X�,�o�+�݋i+J6cZS�
#+�0�\2'�0���%r��y�L�q�}�V��펊T$�Rp.S�Ӻ�'���!j���S6D��n8\��.�M0�!��~һ���8�L��=�i��m��rD�rq��TL)s�&&	�TI�8����4�V�7�U��C�tb�- "]��p�˶�LO5� �������6�^[��&�
�s��g������-�w�֒I��YN��d����9ӣ�h�5�)*Ҷ�\+��nP�B����U��8�;�2���%���q���şK\�r�+�u5�4=��v���oh�)ٸ>����g;��B�m�'>n�_1Y���c�E�T-L#�gbsnZ`6�PJ��֚)H�ƌք���ԛ߽�2�SXE��9�����N��4��ߨ��ng�o����/��%��{����,�qH���\���y����w?�h813�O75d��֍
.�q"8��23B�4Q��<b����0y� ��L�R��AD�h�$�'�$���,	@�ZUT2*0�&��V{t���l� ��~E�~"Uko�S
\6G��F�� 
�����\��Y6|32�����0���X �^P�a����$�0 ��Z0$��ȑ�+��=[�K�'���v,�N�u>����36��*��j�)�2�2�שIa�2/��q(b�� �	׎�U��Q3��4�r��ɡԥ���NA> @�fa�̈�<�^Y����2��j��K�ɧ�ndX�/��3� ��J|����vt}_�4��^x��u��4YO�U[����'���w��B�n���[�-��u��i8�O��t����)$`�������d��|�/���]�o�0�*�e{�e��`x���[��,�%{۹(*�z�<=�d�ĊRi��-����dFO������l���[�)-cy���d��A|hN�!���Zq��Gs���h!}f	ȩ�[�;�^*���q�#��,���~= �Ip]y�t7M�b�.T�q��9�B�r��BU���c8[b��8��^�]Ҁ��S|���T�bBa��ȍ1����/ �5u֤=�(
��k����'ί�Y����{�x��>+҉;� V �znk��'������W����mq�T�
�~��4j4Z���B��M��c�m�w�!J<�sYc#�p%�!���X�'H��'�hP�"Pf��^���%k��Mh�N#����F'<�%!(�K[]�W������T���LV����U!)C����b;�mxHr,t=?(D��0HFi!I��v>2%�g�9^�?H5�pO���[7�3y(ө��Nכ�؏�D��2I�J�0~�тh_'��k[�.�����sC�PEz�
!i�A�|�1n��t�71��8k�W� Q�iwէ�p�XF}����h-F��=0�-�Z�}���S�8�0s�t4IՌע�*T㻪X��J'Y�<"�'#�԰��?o-�XVp!〉�<�~;�
6�`���e��,9��i,�sm��+$ح/�T��܋��*��oW�4��/5y����[�Pv�Z����8�!9Tn)�㺴{��R�,��n�"��v"~ω\u����,ͨ1�N�N�RȜ���)8���bπF,RC��h�J,q����n�Π����N�im6��8��j��-�C��c�0Բ���p��k��hwly��S�6��cb���h��_���l��~�C�6����(�¶� .c�!	.]�?zX���d&�XlxVHYEB     896     280�F�wwa�o��qAHV}i�N�n�x�c�Kd /�����qWv��7ȣ�7��9Uu�>�=�c�]d�t;���_/�`2�i����|R��	%5ږ^&�s�i��u=>;uu��)��Y�CS����S~���S��$���d�:;�e�?AD:+�߯�:�o�E�Rm���$diZ������D�2���^��%�g��-�e��n���p��_��S�gF��O�na`J`J
��\\���~Y��[�4x�Q��z�o�$r�AH�v� �p�b�e˙�2DV�O��>F�A���WZٴq�k
o�M�O��W�po���ؾmG�*,P��\*�Ńz\;>������U]����;�F��g��1T�FO*x?:ڟ���_E��Q�Tn-�?�a�F�BD�}&��W�9�1�l'�-Հm�R9@�lh,pF���S�T�i��~�PԨo���u/}��n��x��a��$����@�l=co~y�j�}���E��G�x'#��y������x��J5�}��ﻭ���ŝ޾�?�d��l#\�{!�3��98fZ��#��a�Dp�؜x����6H���݀�gy4Am��swm�,����K ��JQ}�)߿"�}2