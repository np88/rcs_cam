XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����s��J��@O�L�5sD\��Ӡ^A�(7�8Ax�"�!� -X|�e��������	�ר��A����ݟ[�n}	!�T�x�3u��c���<ƅ����Gt{ˊv�ϧ��hil�qHy3��sov�#n ��@�a��	L��5�C޺�S�Z���GΤXm[��l^e�֊���U�pVӧmB�|�m5�QD��x�Ӟ��m�ʇc4�4Jh�G��b�aHw�3n�,������q��-����z���pU@yh�'}�ܫ�Q�3gU��>yv�y�d��dO���T8�D����B�h���j��X�����rEP�d\����5��o��s��g�Ƚ l�E�1ォ�E�{��_b�?J`<�P��{W���_-_�2��������,�m
oS�v�����q�L�	%Ǳ.��7̱��(�0��H�},�T�'_UR�n�j(<f���8aлy���:���
梶��z�ӻ<J��4J�i�ަ��5hGZ�0��Z�ɪ��d+[:݀�m���m�­S�O��j�Ⱥ���":b����:�.	�g^�"sڴ�?����y�,�`D~&b^ڛ�IP8\��ev"B����j�B��AE8GF:]���o�'#�GB�eua�߂.�]���Y�VT3���l����kS���~���Ϭ2��O�r�cs��s!3��3z��b��J��F:���6�U������{e����U4����
?^U�E���,�6���$$�����P`XlxVHYEB    fa00    2480LUƞB/�5W�u���N^c�S�����G��e6���1W-V�B�%o��X��H�Bax9*K�����M��?�ZKg��/_	[T�~C�q��>�Xqo���y)g�+N�l�QN���Q��2��[K/m_XM�+VW��q���M�OX˅�$�a3K��V3u�.�xHo�����0����Q��vNN�sv*B|#� ��J`]=�Ŋ�3a�7���z�#j��$*<lە�9�e�S.#��"*�;�-�2�a�\\P�Z��b��F;k�p����(�0��=��-���
��cp�[�j~��>������M�0��A/����Z���v�>-�v�yE�����}��B|qT��[ކ��\YL���I�b|�p�8�3^"�A�V�N��8A��Z%~ �/�{�E�al!�����m͑W�\��V̕�������d Ʈ�B��:�0�(���\,��/�94�C��)N �q
��ɳ���m��$��8�;1�G�pyN�(\R��Թ��	�� �z�S�%8�F��2�	kLoԲ��辮]�s�����8�?)���C���a�yƖ�Zk�rſ�w�38W�������
�}�9�K�@���ѓ�X�o��
�x$�	{i��m���ֵ��w�������LQ��_|1-?0_�w�j���[�W%�㵒ş�4�~���
��ƭU����&F�u�[�~��_�A��ߺ+��-��]�7�Ɇ�����x�&�!1V�~3�-@��|]I��E��`'�{�l��~^<5�ú9�"����?ud-��ݰ��M�H�`���I��# L�!���vÌ�X@�i� ������Ji���i��n���D ��"h��8m"ȌXDn4�<��v�	E�V0��ù�L`��b��Ϋ���c��Kh�ΰP4@���O���ړ"E�g���� �Ǡ<d2w~&�9뉨�m _ػ�aI"9<��� i��uD�6�Y��b�2_��o("R�2�RQ�e�A�y7uޢ�|�i[���Xy0=YY�x�H@y�1������YC��y8z��T����[��Ǳ�H0�� '��������JRP�M��+�K/��\݃��I��۞�A4��W{AqWؔ�z)�B�^zT\ȴ8�� �[G\�ߑȗ�oi�@�A!l���Ɩ�
�����B��M
EK�gTx]Mdf]��q�:�xoC4��6�<FH'C�ωa�F3ν���K��8��P��q^;�9_b6D�3���Eg帥/U�z��Bϸ#	pH"�NR�VP�άLB�������}%�_�����Ha����
Ss7h��NQ�V;��wE��lA.s�{r7j6.W/��6�kǝ
9d�J:�${�S���'#�r��Ce��"�4���
}|�(���%T���@��!�� ����lA6?��8b�1>���*EL����$�+Xfv��1����=��t�<�ě�g��Q&�����%��W��)�����a�8��y#�����̵vOZ=�)�2}O(����4ܽ�(�����3m�2|	��n��/<�r�mT��(M���u񸏧�`+�'��v0U��7�dt�c��#گ��V �Zp�!t���EO�+��W��=���qrd�:�s�#;(�ޗ�-J #P\���"7��^-�;�������٨0���4�ַ���Eh/�%(U������w¢	q����[n(H���y�,F�05�7��_P�K~��6�-*�e�-x$|�g��X6X(��B�%Sd�6�ҍj�����jĄ����!��pM�H���Cȅ\s<u��gH �#~�q�
��
<a��*Ib��ǯ��Z�K�c��Hz��X1�;:���V�[���|$�L�a�Q������I6���^hA�ҥ�"%��`}���Ym�,�*�U��<�,��H <�|]��������O�#�FywyvG��H��
+�(�+t���7���I��~����uw����ˣ �q�cԴ����юʗ��?Ϗ3ǺR����8ڧ1[g�2��B`�,�۫7��vW�rvi��ф����Ӝ ��\*�� ������0�dP�¯��g	�h20�[>X_�4���d_��,�Y�*Զ#F�*�����'8M!�[ՙ�7���>����+��Y���Y~�'<v�%�ҥ��i�����L�`��j��.w��O-}P�N\-L�${]n�_�݋�*��(۞��#�$h�;�6�ლ+�C
�1��"e�a�2�6�
�]S�u�.�K�C�Z��'�([�ofu�m	�`E��]���� �#~fƱ(�o� e2 �r�	T͟B��y�ΙC��Y�)I�Hq�LM��!e�,���ǩ�%���\DF-�j�zM'a��:J���׮�1��Be���9v����Dvp/ȱ+�v���I$�L9��@�RÚ#�9@d�����&�2}��W+����̦�l�l.��EO�n ����j0�;oCJk��Ox�D�C)-�9˘�U-1<n�M\:�2�Ѧ樌��񷠫�'?_d�u<&w���#.z�'�?�:���tc��\����q�ߋi��7G���^��f�xR>�.'��؋�z��33�JJ�M)!��؊�ki"b/�����X_l�x��X?u_TM0{59\㑦�d�=��`/}!^ƙtþ�N�~�꽛�&9i�V%l�9Pq���Zg �V���3���}�ŭ^[�z�v�P�۶ y���D�124͊aV��E�C��bQ2��И v�	M�īE����w,�D�ķv������k6�fP��Xye���KH~�n�)�;���M��P���W�qǓ|Kq�t�럦4��[���j�K�OP�}����e��C�/p�tJ?>�HT�nAA���Nw��o� _�߭����D]������5.�5�h �����^�d�ύ��*L�?[�<T�۲���a(`{π=�)�[�'��m��n�3Fet���xO��MP��n1yjٴ\�������,��ģ�ah�g�h������B����㺭����rs���q/E��D>��]f�µb^nOܑHh��!S���'���]��*E�V<]hҁ66*�DG���W舟:�g��㤏�sG�h����>RG��$ov�HԱw
ԨKٟ��o�t���Q��G�%��?p��O�^�P����氂m���9����d`�P��J ��{��vbU����K��ue�W�����=\i*�{܄���'�J����+8�r}Z��oA�1����u���ڄ���qq�,F���u%ә՝����0�o�����+#$zy(	�>�M�QYd\���w��\n�HjV/qԷY�@��x묿�$Od���ܨ_���J!,��?A�O���5�|0�ڴ6�_m4۪8�(��dk��0�db��4���U�^�	�ZJ %N�͙�@� X�u~	0ƻ���M���)�JLȫ�y�I���r������J�w�P�鑜Ԕw��2���DW�/N�[���5�'�;�k�H} sV�r|���0�h<�[����o:#,�1��ULj��gk��k�	�@
��B�5]x8ڙ+�IN�=Wo驇D��s\���4��?.��;fD������G�$��#�iZM�

��k�NT*w��Nm��/�W h�a���`_b����{FK(Π�<Xf`�g���Oc�B>r�X��vl5B3����jV��@��Gw~�&9�͓�s���(�T+98)_�8�{�U@B�k�����F�\sfQ��~��/b߾CY�ܯ�e�G��#%���qY(x���v0��J��T����Ho��qu�:��(�GU��i��/� az�I"_2���1��%?�s���B�q|���ھ�5�u�L�Pn�]�[^|� �)q��z<��-`�~��S�~j����%�7h�@Ur�)E_+|���tۅx�9��z����Ǳ=-�6��p��;�7�o�e���2�+]R�p*6��	(e�OH�	�1�̷F��[+�3�I���d��Xg�e�W�I �3b�4���Cc��"8cΣ1��v�Rժ T;AHe��p�t
�(|v�����d�?Պ3��fю^�^'sF��uۙ�R*�v��	�]��V9� d�bs���} .sб+i ���ٸJ* �WPO��G�!��m�70ɣl�&w;� ���N�¤Y3��m�5���[�=уs�;�s��lW�p)<��q��Q�:^�*3�-Ce)����Q��Ms�V(�:[y�D˂��J�o/NC����f=R0s�������W\�N�
jx;�w���;j��hɽ���b�]}a����!��tLN{�������h&䠴�U��R�^T��7e�#�R6K���:�����ʬ8� qH�P����sK3p���B��~�W�	U����(�,Ts�u��J"���<���*���/�-�/!I[�����5<+7��Ln)D��r��8 �cy��E���5݄�����t��mႣ&y�n���>��O����g����DeO|�Js����� 2|��T��X-[m���6��B&*�����3.�H�fX����Wc	���t����O+3�+��S�-�,����d��[��5�y����5�p}@�G����%�<L�J{�~.�8�K^	l鋼��P���%�k��VRs��1�Qpid���]yAJ^�VWF��b��X���<�?.��!?2ѯ�ۙȳ���H�����7~�˵~cA�,��م$tY�KtO����=iQ��܊K0~9�ul^��V���A9̚�j̌?
k�pQX�SV��,r6��B#�C|��ݿϖ�M���3l���]�#��|�k��jz��I"�0p<��zX���0'W�q���ɸ�3�c9&�����]���O�-��!�{�M������W}��+[uOŮ�(5K��m�<1��]��rv��ya�ǌ��2x;<���r�-���:T䴛�0`�50£y���è�����/T�寤0�>��ie���V643"9D2��m���d����&ĩ�rc����7^�T��Y�����P�I�y�'�o%.k}*8�0�B��g�m
_�A�'a1c@&���+��R	�ј���%�ƌ��f�a��L/�G�z������`���3.y#Q=B݂���D�;IOOI���k���E�"f:��Eȵ�:�'ȟI�w��#֛��gI�pR�>]ye��L���q./pOp�T�"�?ͽ��mW��r�o�s�k	�ۄ݅ �l�I�x��J)]v^~�<:E'f�P�M�G�\�t��R� 8��B쪋S\�NpƊ��? B�/�ϙ����,�P<���B8&�d�hQ���3�PR�� ���X�n~߹d���6�a`g֗/B��P�k�74��K�os���]a*#G�(�Y�x9�r��f��g)���@���mp��&�b���W��2�_��&H/��w?�s/A�����&�F�T�]Bus��� �d�s��@س��o +��2��qw��
y���!~f�3y�t5���M8/��ąo��g�\�?`���M�۲F<�ei�A�9ӓ�d�7
����d3�R>"���~�NW�`VM2d�~�� � ��6;�|=kB��S�o+�A2\�����ێ��R���P�ݵh�,��xu��o?J�ϔ	6v���~���;��� 1�Ji�Û՛l���E���#���ѐC4p�H��[�Rk���K�b�1������"�����
���Pw�\�w*�V���N�U鱵��IA�U�p%���o�V���V��/@�tzOT�ȩpLn�����GQX����k�mԶ,�V_�.uv�'D���[�	Q��xQX�e/I�x�z2	Mn0�����.Gh��q��A:�|>�%���bmP�7K �P�L� .l��Ո��n$x��C�F'a-dd�.�*�I�O�8i�in�$�i�P�굪��
��tTNeh��&�ZHMxw�����G�G�뜦s%}�ܧ�����\�+��׋��M�b�Ů&��?���5Ҳ���ܶ�N�H�}�$v� �*`i!U��(ƹѱ�0��E�U�%�:�s0ߣrC��� �jsь��ŋ���F��!l���)�[����d@�En)�L��PQ�������`�vYZ�v��F��Zˮ�"�%�4N��Ox�l�%�� %�3fH��-7�1�I���v�ٖ��
5�Ş��<��M@��_<�Vf2gI�e\��o	k`������Ƙq���!��+�km4��M��r�LA���ʨU�8�n�O�%�����䪖�"D:)�v�F�q�d��~�>�GΑ&`���M��9D�af�D4?EO��h�*X����<�bmެ�H�"Y���H�����V�Owc�l`s����~�e�Iy}�/�&�7�O~�bH�s�_g{���~�U���c�|���k�ׂ���-)��)���ϼ�F2���3��A!��O{[��p���+��m.�c�M(D� ��v��ʜ��0#�@BP�{P�LlW3d&Μ�4t��KWjl��l�!�Wϣs�k9��Ĕp����o*�)`��_��Ou�R!�+6�lC�"�C�����qr�U�яO�P5���n"���'���f��[�o�Hf˯'"�O���f��9u%���1+,?nߘ��FW���*|�Ǔ�Y�0�b��-K<-.ޑ��t���]�ܓ,�e��*Qos��1��㇏�No�Z��~�w�n�*�(j�"A�v1Q)0�_r��.�S@��Y�%h��!2jX��i�T%OrT�Tpfa-�4�d�� ɮ���
�y��TL��{�}KAU%~���<3���I��30��&��+h�oH)�ܩW;_&�O�e�+��9r/cDX�.Ӥ�]��\?p����g���%�Q.�����!6�mx§��"8SR��2ۇ�el-6��Ara����3�*���L*�;Ec&dff�TCXg���!����%��c4jl�B]ؖj�T�!����+:50<O�8v��:�s)Օ��W�p����i��]�~����k_�OC������4�2��^ݶ �@3:̻�g���ƶ���fi�C w���R���Z,j����ސx�P�U����/ ���e�䂧���eӨ���<�JT�Q%ͦ�֣��8e��`ᛊ��8RWZu�$D��ۉ`�ؐ7F)C���%v�Hi�6ȊW
�J������"D���]f��|��e���_��J���~5^��mv6�zЗ�O��U\��@��v|��\�K38���?M��r��	����ȷ��1�+�d�:����{��y�ŏ��#��,�1�7
E751@�1�3]� ���-�&��8��۠ؿ.fM�Aw>��Vr0�P|�h�4�d
�)��CLѧT�n0�a�����AmZN�E���Ւ��{��E�3���|-���}����ń9fi�G�s�S�T٨�ծo;��8G�b��M�d��w�����ϛ�����?��L�8)���)����MI\M��WD2���	�6!=���f���t��^��"S�r�p)П0F��������0i:Ĩ����G��jY<�kD��s�O�#+f%��;����0�֜k�W({��X��$�.�I����6�T}%�^uO��XMK�<���<�k:���D_�7��� /�l�n���.�3�q��ʴ?�ArOQ�)?o���k�.!ة��	�o�v�Ց�-[2սN`)Mhr���=���(Z�YP��WI�wbL;���]w����W�tJM�߾�q
d���10@�MJ��P���Tp�L�e��ݍ��b�V�|	�gaH���k-dᅗ[Ƿjڮ@�ϿZ '����o�:z�V�Z�n9]^@�?X.�*'�L{/��H���pFIU焙���hOm�#|V���v��+�bsCx��ϲ�i]KG�(�����kB��yN;F��( �`�_�uD�@�av�琬ҙ����l~�.�Ȅ���^�L�&,�E Ϧ}�&G]݂mh��1p;�QXec8�3gP�^Hjn �& �7Yn*ĭ���V^C�� ���4̋ea��O�����ZV@ ��nHAk%4�e��m��ذ�R����ȣ�ͦ�]�+���o�z����m�m�rV2���H���X{�ČS�AX�ݺo	�� U��#u�y��ŉ07Eٚ��������-sO��(�a#n���4Z�C8J�e�%"���Wyۧ����.w�ӽ�9qEUF�­o�1:Nєt���$��ߏ�Ӣ��GEܮ��UH
�'���ߑ1����F�u����,������.��K`��ZHu�4d�(:��3�{ZPKFMJA�c�hp0ľQb�㻉��O	�B��ٓ�$�;4�$oz^���h�Π?�" ���9�+j}�rST�8{�*�:i�mg
���z�( �o�w��rU�Xq�Sd�~~w`?�� ��zM>��2��^J�ջT�
n�-F�~�k|�@��> 0=ЧY�9f�X�"c�5ϳ;�$�_��d��V�)>��+�a�2(%�O�V ̬�W��k�S��drR����!s��Cv�Ka�Z���_B�i�C�ޙ[R3��X���8;>��I^���B0e�5��W{�=��
^b@�[R� .�`f����pU�Z�`Q��U�楯T2x��ُ��fL'>�'":��*���$�w�����Y6��&_$���@"��	-o��;��A���A��i$����?n���O�T�t%a�8�S� �	�ͮ�M���5z�`�"�UT󑶛�UC�`M�b��5�5�R���M�7K��xm��M}�>�����Q���:tت��H7�{2ϫ������Άr�]! e<8��'?�⠛��١�q�_�1�7�f/�����;E��K���$ư��1,Ŋ���X⍡��jK�g��:N멵K�|����b?C����`�'��Ta�j�i�d���揅nsx�Ї�t;.�v��Sڽ^q�Zp��s����缏�ۈJ��x_`q�����&9Û��$���e�:��0��t={�_�7��	��l�"�U�2�b��>i��v�C��蕬��QZ�CD��]����x,6 G[j怪�wc�Ɠ��H�2ټ���(P��k�ZV�<�4�(����~5�Mo�K+�R�&v��z��XlxVHYEB    964e    1150�N�Ԋ%����.��8.*[�N3F~�	O����v������$$�æ-�ڲZ�����?�P���"�1)Ke)�@����y���ז/]�������a[v�)�ꘕ��gN#���T����u6���t��վ�������i��BJ�wS�D��w���r\��D�2W�(I.뎃=6������f�d�ğ��ӓˉ�s�jDm9Lmc�;����̃�E��z,��fB]�=�!A`�Z'��� ���crQ��3�r�4��kNZ-�͡��S:�_;��B|�|2��%�����]g�������E�]���ZBъ@�� u���M���_���:<�4���1�-�cz�CV��C���ZW��0� �Y� �>׆>k�z���=�
�J:�L�Kp����QP%ﷱ��^M�Q.���H�N�9�`ƥ�!�o�h�
nh.u�@� ��ҏ�Gqq<}�$�z�y i�?�Z75V��f�'�L��8r��m=��,�=�y�9��/7#($�6���zo�!o��"0�6����u�gp(&��ڊj)��Nټ6?JA�g��9P�\���&]�KI&��"5����]���_x�+�!��7zf2��.�FL4�q����w��S7�$<�� W����؎�~�#�P>E���]>9`��y��r����UV�lP�����u�V*�R��������<΂@����ݞ�u�MW��OK-��Y�7�&W�uH
��S2�oZ��$���}��,���,wSX�ޯ�,�`�~;���|%��%��.��"�S�������E{���۶ݸ���ܐ?�K߿J@3�ѣb՞�J�^���N+��;��qŗn�nC;�h���Ju0�̀��<Y��}�7��_���P�kt���I#��X� ;�Yέ޺�W�z���(!>���;ӡ}[�-4��CR���ǟh���w��ih�R}���J�I����w���8fgq��/�O0��@�A	�a�>�!"o{� 'Ո��� �u����u�-�q/��kϮ^%� qV8`��v�B{�N m�;��7mnΠ�i��T'��¢f�䛴�VÑ߬�>�X5[K8.	z��X����oę/X.���S��`�˔���
r7?�
�,�X�
��1�zq(������#��1	��wB%��Y�o(t̮�	ϝ�ћ����'��˒]��K$�ub��D+�	��?�_��`$��XO�����ҍ!�ۚ]3�n�?/z��rY�*��zLv�mG��#/�˭p���tc)�n�V�i� JkѦ�bz>Y�i��.���jR���'S녌[�ئ�ZGh�0���-��N)=�ճ��ac��{��T�����<�� $c�'&�0���%m1Z�Y�+��Q�f�$�e�u�6��k�p��Cv�Q~��S�W��Dx���Du��}�6��8�����~�d��6^*!�u�h=�޴v%l�p�t�K/�:g�}�d7>�
Xw	�L�e��6��DC\/��GE'�=��o߳T�R-�M���oA#��j��	��	L�		Ә}�auiJb�W��3���v6F���6��!W]�m�A9�
���O�#��/$�?�+"���M'-����]���t�b��f�+`:�a����^4yB����!_���@�?X :؛؄Vl�ﵵ�\�Z��0��`��d2��cV�	(�R��#P]0���mm~0a�GفW�N
�%�$A�{H�T#:?������\O�5�����.!����QD�1��)w�}�{����7:�
|\�b��ݖ1��&盉[h�#{��|�HԴ�����)��_�L2�gS>#��x�EW)`�s��	��~�@����[��\^�*p��t`Di��%���,+̖�����j[X�q�f�:�rY�m��u�l]��{cZ���?Q��I	,�������w���B���e��g��%�;kTR�"	;��	���h�.:�Z�P<����Β�-���/�A�0�H\�tr@V�k_���+��ہ�n���m�c�۞O'������L~��=A�Z�X���l�p\�4����;��u^ip�96q)�R)�3Ā%�%ɈAv�l6*&K=���'$��8��iF�;�^�m����C�f��dS���6e6�B�����ta� $��	Q�!����%o��ה
d\�����q�r��LlME.��o��^T�����t�y�����3P��ZV�Ưk{k%�S�.�$^S�%IhZ��<	P�����\��Z�S\��� ���^D�q���1��J�^s�uL�����D#kA�q��²�kg�<���A$.�;�;�p��u��uG��Ut��LW*�I%�[I��(ccs� ���8Gѐ3~�s��38�E����/�B��i]/�1+���B�R��9�F�C��|�����_���9Է��6_^������Y�[Sk]<������Q\��G�Sl ��vg.��VƁ�zUU���Wو�)�ʸ�AxA��I������פ��T�C4�������1�.	<��t��v���U���y�1hfN�O�6�ޚ�$&p�oƤ�X�}�j�������֤q��0�	gl�2D[�|�"��сt������1N��fߩ/s�V�?"�~*i�l:?�Q�����y�Y�*���q�SpSV�9X�$�;��'�j��Z¿v���ud��Gs[J!�鮯�i`�$��Ǿf |7���p�f~�}�4�S&��XLd�uӮ ��t�$�������g��+7Lל�UEC�0�?(�?9�9��`&�����˸V2SSc��$6�"҇����lM25�m��@��$�(|�L��`�q�T�_���H�z��n�@�Qr�-ԉͯn������7>ɧ.��#��!D���
 U�q7 ,G%���E&��p��Q-4��
�:J�'�Vp�U��ْ����m܍����ݿ��*{�uCޭqb�J0<�A~Z^��і�^濏�I���lĎ�"�9ų:.���=On{�U�S<�]Nid�;R��y�D1����9���.�߬6�|���y��W�m�?�!
1u�M6J�u�~Mޛ��:��Um�;��:?ʹ�r�w�Ԝ�S�I���
�FF�b��o��bZZ �L�;���Tv�y�aC���;$�_܉mϙ����xϹ�я�^�Mo�z�}�o��P=0p��$F��pY����+���f�4)�n���8�U���I�$��"��FQ>�`~(�	aZr'�`�������L��F��d�x	w`N�IH�/ڟ_��_b��k��),0���Q��	�mc��M����D�QcH��-�i�?|hO��M�ka�Џ6�
)k�� �y{���BxU��r*Z�D�Ğ]��	~�"h"���c�O{��Zx���O��jg$��RElW���}<�_�D{1�dO�t&q]�F2�>[�x�N�	�q�`g���/�("�9;�A{�-��0��s�v�o��*��`R��=~+M�o�A4ʫ�4�#�6��W_���s��q>ޣ�\�֨�;j����9�b7~�;����p �R�O��`�{5�J� �(�8~s��ϘA ]%��
-���f�F�c`��w}<���߀s�*�;�u��ES)^b#� �M������g���r�V����[���(��!fuM��8$\�F&�v��UIe�"=\�������n�A���p4I��Bƺ�"o�0�Φ�	IaX�s�!�ŨG�!��@�8����~+�B���ޘ����X-�v��.K+�)����_u���a��@�};q"la�VY���j�u���O���Ej_	���e��R��j4f����\���^T)��[(`����ܒM nwh5�2���.Zc��Uc�� ���/s�w5Ȏ�V�������7G
�e>�m�O��ϙmR��Q�������Dn�<���}h�v�R����_���]��to+��gY�,���EJJBw�BX��㟄r%Ͽ�N.aJ79'�N#��5Q����myAf|����>�ӕ;��������;��6����m�/�^>��s
D�`$���`єdȳ:Y���k�	��0$yv��w���O�'�����|h���p�2Ӈ��*U����j��(0��|��	��ʘ�O��mܑ ��v�@�%W��YQ[�L�<[k�������V.,z�zT�/'&���YRu���/���[ء׌���Y����FSs�_��R���&j����d�$�k}��vIB�#{�dF�`���+`̷G�0t"��Љ��Y���9�8