XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���Hs�)��p�"�t�}jZ�����#W�K^T�2�u̴����Fe}i*�7��ͭ!�*x�ʯ����*�'�0����!~�[Y 6��}������s�M��"�������d�6f�Ψ&�.���)��{عX�蹣��Y�qQ=V1�!����2b���p��b
K:��
�ܛ�h���^�vf�I�ыK/�z�����;�paEKW���F�Cܐ���JE6�o�oa�Q��yJ��M�.�S�7G�dv���|�rl,�&��䮨B�.��Cu�I��G��q�&`������[
VzmN��^:�ʃt������IO����}�_c��7�2�^K��n�2��ָ��ϭP�<���hN�nF��uX�[���-�)e�Q�8m���A�W��M�~Zfn]aݼ[%"�!o�uA�3��Ҳ�T��{D��f��M�G*�_����c���-Dv$t�>_��8x &�`UtR7N�-��F��Fߒ��	��ܕ Z/t��0���� Y�y��zܞy-�1 <Pѡ���Q���W�F�vG��$����S��^щs��xI�߿`�P*?@���1@V�!wk�:��'��� c�7��s�Ǆ�z��������$%Qc��5���{�?���@
����蠥@�����kӠ�I ��X�q-�'��YO�6tV�Ʌ`����M��^�0D_�)��VѠ�����Ie�)�2PR٘�[3mk�������/��/FXlxVHYEB    fa00    1f70�@<�7���d��_`(U'G�XO��"��Dؕ�E��ڦ�ݕ��!���Ȫ�A����F�:^����pH:�����ӷ��76]^y����s��Q�P�b�V`I�"�AU"�2!�O�g������4���%�`IbU�^��w�вGwy;Գ��7�2�lK��["V��l0#�/�lPb?m�1�Y9�8���%����!4�@f�YƓ-H^��#�1����򪜕{uA�"B��A8T������n�P���N�՝gS����5�O'_F_R�1i6z-�8c+܏�%*Dgu�i�ϳp�"���W�!�]n�Ĥlɘy�#L�G}Mx#��k���B*���zN1�J1�Bx��G�PV\�o`����vx�2]�ji�j����$�2�� �S1\۸ <4̽�"�˖L��j"a��z��ē�5�j�R~�	l�l��b�L���Z�W:1�����oRC�l�gg��P,�,h��tt��?��'��q��S�ȑL�fvF������iN����("��n�"��KQ�*����LqG���' a����x�>���Ѽ3�����h_�m��fǊ��q�F`C̏uRD���dJ2;�'��R=���z�� j@L��/W�H ɱ��n�Ÿ�D^���ǆ`?�i7�����R�v�X���A�k�)T�Έ0p�'���V������c����M}���b�m�Qd���H1��fR$^���u��lEOJ���U�֑h�5<�&�ons�l�"�F=��.hpĢ�����PP����}<6� ��-�^��F��چ �_@�Wr��k?�_�짗��� ~�xpT7���S%6�i-��!a:Gg�RIx��N��b�`\
�5edb�;Q�C����b	�� �04����v�a�{QR� ��M~N�Q�=�V���51|�d�h'U��s<���.E�=��*҈����TnxN˒�D�G<^ō�$�C�u�"Ő���k�Y���U1��Z��m �+�+%�|�2f%��S�i"�m����#�'f%���L��2���K�(�Pp/+'���q�����鄝���E\Pl�>[�~M��`��h�ԏ\X�o��YX�@�๋/v�D���˫1����3j]+B��QC\��g��s���?hB?K��T{���(�x�;0��ݸNPF.=��x�S���� 9�/���%���ϗ���8S�l�s]�0�^C"��3��vO.8����	.��g��������ZD�U�0�;�7̕Rh�@h6rb��};�y����ղ|u��)�����(K���uE��,Į�;�jQP�B(z;�O[j�	,3��>>M~~��ډ��4L1�k�b����T��2�ܯ[�;�R�\٪�<fX���Q*j>Q-�7��7xqV
�i���T�U�/dM�RDWO6"��m~���F�GQP��Rg2*�a'�y�c-�%�0\�r�T~�j���{2��(^}9"_F�Uyl������0���Ϭ���ljͫ�Br��h������w"eX�v� b���`�ߙ��`Tr<�C��('c�d`�)h�:�+��T�̾5?�Ł͂i�}6�0����Rjr�벟��R�\Jc|^8Q��x�ٮ,���ʅ��>�T���+y���ĥ���s!$��g��i�y4_�(ѿ<�ym��:$�l�E���O�5"C,pp�ڇK��2�F2�Q68�\y)�H���YDh�7��BF�ߏߒ�i��"~��o5��=2,�s}�0���X7-����c��lo9E�(�8�E���@�I}gR��B���h����mǏ7E $�N���q��n��B�D-3�8�����o�ܩ�8�|=j����6 GH�����u���8t�͓P�v�xT3�߅�1:�%�����������S�Iɽ��ŭ����7�nZb��i���~���0��2P�a�.�@m�غ�uς7I�5��01�@&�(�OX���Y������6�ts	u�^I���W��Y�K�s���*vPs�(o����VN2=8�FږK���E��}c��l!N�^��7���M��<��{G�/��gs��Jԁ~fW�ð���j!����"�g�[[>2��+�6�����bVє�?^�w鈴x��Qߵ��1����S��>���0���7��Ι�9h� ���^�?�deذal�lQ��)J#	׈#`u��������v�I�=�4�(q��jGȃ���,�;t&KN̂�D��3��p%on!E�2%���Sro��.a$�����N"`�H�I�>�b:fm�4���ڡ��ղ��9Q���v縨	�ѕ�MqGC�$s$T�xa�x��C�>����Z����L���ീ~DwM$=�A��0z�O0�>Ge*h!Գ�����;��У8�͈Y�o�B����̎�;�m2���A�3G[���:S5���,��B�[e��y��ڷ���X,�Jj���IU���)[�	�Ycn�iϐJEq�f g>�ݒ	�k�hV%fHI���r>� �Jya&/"8�e�N4�h���s�I��ݘΞ�綬������p�`(y>+z�d�y���X�B]æj�c�'5������A;��`Y|W8	�-�[8I1�4pYC��h�Ow^�9���ť�BD�f�9�r��ٮ�f"��/Ka���9��#y���,�/q�9�n� �v([�_U|d��W� ���Ìlȹ�vYG�3����dtt�:���=a�jc�6s)�GV'ϋ?RơȨ�+��sOr�$���*�溺�D���0L��-���	���_^��a��kfyHF|�����ر��N��=��g��S@�z�w)�;ȧ��v��Js��yo���.�*a?�/�@���=�v�X$���Z0	���O��;!�!���G,�)��a`#�x���q��c�:�e�'F4�_�`��m�py%+��j�م��������\���!�8=J���7��jp[5{�}j�@·K2�����ܻ�ۏS�p���Ռy����k�^��>UC��f��?�քk���X�~
�m�.=���[����Ӌ\(���R�.]c�ьU_-$}�m�[@�����`*$:4X�{A�?x����1�`nӨ�ճ��oRJ=�W@�sq?,��d%�1S�����(P8�hD�A&�c#{R!��l6�6�vKߠ�=Z�4��-1 +,C<��Sa|���W8���V5^|"���NN��qgG[�C;l�	��<~��B�� -��Ұ|�!�S40�v��U��CKG���2��jd�x�g9�k
J2{��K��!\(>Z5&ڠnz�dy�T㯪�0Q�W��E��t�y�44�5v�CS��7�^�*"TI��mI����cn���z3`�����-L�������AC�\�yݺ=��S�+Y����鞴�~��i�6i����ݴǩ��
��h&%~�R���d���/@l�~;�8"�u�7��x�pA��L�Ȉ$��*���>.XJr��.�n����1�a}����n6�m��bA�mY[��\�m�n�܌m�{����wu?@�W��-�qS궏��H���kta��<�ں�<s�Q�o��<���� f�&HYz+��Xq�s������0�  {��1�j"(�O/�%������i�{��R�-�����I'&�E���0I��iHl1���/��Э���=�_ƕAJ$��� ���:��g/T�JϑK98�v{��:�*�i�>2E4Q���S� P�9�ES�s����H�#v{h�Zgqh7���)�`�6�{�A����5P��ZY���P'�+�'y����B��B�Z2iC5k�W�L�>������.�h��u���g�C%U��^��;�8���fp���~�u)[M'8 H��_��b�@76�f�a�<�k�H̢��^\��h�Z5��9�Z݈��`��q�"a�YT}r�>�o^���-k��͜Z��<R�h���x=&	���ԒZFg'�A+v����Іt��������E�yKL���=�G�MV�[uj����̠�-8V®(�"�zgZĊ�ǭGE�6͙:;��V���o��Ua�E��qS	�����1���0�tX��*��_�m>��Y�Czo��)l�'g�|_��}�!E.�/q�NubW���7��h��0
�v��,\;��H��!v�׿�d� �ěvH��/@���Gs��B>5ā7�V��URޠƛ\:T�	��]<��pɍ՛�fq�[���͜����"�СG��)V.��C��dQΥ�,"���',�h��y�J��EAȦP��n�tG=���r�T�lE�{d�MN��䉫�C�[���W��b1 N���+'ˬ�̗`D�4R�C�w�=��,�;Z�R�ִq("��*�Sʣ��뭌�ZJ/��_n���Ƣ��l�VN煡�(p�؀��&І��@��Tp�Sc��4˻c���7�+n��Cƥ@u�֪W@AE=뗪Հf�:ʕ!|��t�9���/Y�`!���`�c� ��g�a6�����sy n���m���3�9߶��-��K�W�\�Db	P1q����U��*[b݈VI7(t}j]�=�|gyT��Q�J��a�y=����i��~�bmRp��\��Jq����dA?�.��5Ov�$�'/6BV	����B��s��"�5�ѓH�7�$�)��ƚ�E$ᨚ�j$�����~�(k�-�`%��X�C_X�*!OwE%Y�#8A�N'U�ꡙC�;��MxW�ߚ�p�;]JU~�YO�퐸p�05���ʛ���neN�.(J���	�da����G�̓l�Ow�`�T�L���=��M�[������W!su�O�[�0Oo���
cJ��ыPo�%w�(rW�=\�cJ���sD}{��Fl����@&�4��0*�ڬ�0��y�(�v?��g\d� �u�V�So��K�>����|4�I1w�S���,�D�k
[#�ˋՉC����0�iM|	|��5�c��#� 8���Dh e&���Ќ׀�0��]81Y��W�����rjo�����'u�i3e�!��ua�'���a�}b7謁T�t��yn#��p ��?K��3���h���h�^â�$(݄���~Bۢ/�E��S�͘ZA7����]k�R�7㪞<}�������B�7��FQ�g�'��Y���@v��Q�=�w�R��:��L�g���	ܯ|Ф�򩁊�&fD�n:*�=Px�Q�l�}�DT$�ZP��)������aG�&^yJM����r=�#D�x�����]��Am�Ƒ���b�������p�_�Qq��K�!s�������\K�8A�^�L0��p���-���zX����Hk����`�q��{/����&)�3@�IgT2�3u�h���������wV�*��Q�u�b�aY�����{Q�1��% i��q�}���� о�#�F!���uܦ���9h��T�s��n�����u�m�R�Mڌ?Y��A޴�5+4�y�Z���">�xd.�M�1��m��]�$D�����!8o Wi��H���D�H�DJ$�
b�;�i�V]���8����2�ZwɅ;3��Q��.+Īhqx��2�m��ٹ��U$t�F$O|��v�'㉠Iw�!P$�]��c�"c��D�0!OyⳈ]���|C,�fB�Z�5/������a��#����x6e)V?�L<��y��	RQ�ZAY��Gg��Ќ�lL�(�d2JS,��3G�o0�q���QԵ4bE˿Tr�?�	.��@{��6ˁKSf�o���V~)��|�GxYv'X�g�� �#6�'4~j����\bU|�߻}���0&̛e��C��ٴo�|�c���i�����q�o�y�&��د���ǡx�ݽ��@P6յ0t�FI����j1�}<�2�c�N�����՛v�0�9�y���Yvv@M`�`����� ���G�g`[hr[Pl��f}�=j30}",p`X����%��ɕ�m���LÕ,�0ο/,h���Tt�QP��K��3=�����[�S�Y�s\cH����0W9tӣ�^k����.��B�q��zϺS
s��UI�	�2 �B����,h���ّ�=k8_�k�K;0mO.kf;xk��ט��j�ѝ��:��mr����Y9"A\O� e�_Kw��i�f�;�?�p$���I�ơ���B]~�S53�1���y������,�@���$b��]�"0�G
Ȳ�)���3p�ᩫS�8ٻ���Z�ȧ=�HR�̼sv����S ;롞[^Źf�g0g�G�!�o���:N�L�n�>U������D9]X^A��� |<50�JR՚Y��NK�Q(��&�z��Y�t�'�����|_��(!��Q[ɝtgi4"c����8��b��ߍ;w��>���=��/\#[q�dh8���r���'��%����'ڇYL;���N�8���B�����j��"˻�Ԗ�P�"Q�umK��3m�^a!F��H_@�Y���7� ,t]��ѩ���Ѡ�����9�c�{�v��6�)�v�s#f���5ωcr��_�oӢc�A��sz���A MUh��J5��!k�_��$�AK�K���Q�g�2�w!?��3���x�%��Io=�U�4�)X)h6̊�R���u���\�7q��2%���I<*Z��F�v�G;<�Y�>E��	EEt�ۥ�H��%�9���C�`�*�\�%�%�o�5����G����!�#Kn���Y�;{j�R$��MX�Bq_�ƍp�;���R����4)��3GE�r��<���݈:�NP�`�p�,i��]�ۈ�P��ݞ��ϝ� 6TY�vm�l‍#莯�`33?3� -9��fK��^��9�o��nKi�����q�q�Mj��!�o��4��0.��h]��,�!d�Ǽ��;�at�������1�,su��,��Щ����za�N�m�-z64<� �8�$�$��+b�22;qV���V�N<���mPd�~UX%݊I�<�� ���AHⰎ�i�b�4L;ы���5-bZ�!�"F0a��֞�EvK�o�Y�n��~D�yk���AYaL|�%��^Oe�%���9�!��@��K�c��UdR0y�����Z9{���ȼ�?��6��R9v�
��8� ;�����rsv�䍻�QK��%��pn�O�d��GO��	t@����0o��?T�n���U�{�B�Y�PMEn_n!EF�_�ٛ�����ܰ�U�\�� �*pw�<)܋�����<�6�
�OG3-7�l ,��[�Ki2����g ��y���D�^�(�"��ެ_v�����c�%��6,�a�q8�n�Z�	J�y���7�
����q��^]��Q#���:	���|qC�=��H��p���n�
:�qE���5�_�qF��d� ���rá"�|t����:�C��?��Z��w/�a���:��bf��
�焙�[��~G����k�P�<F�)x����|tP����
��J��V6^�UJ�ص���j�+l��fҮˉ6��^��^gE������Ӑ�m�F�*�H��}B�x���W�Q#����K�a�&;bD�hp��#S�H2ș�\�صg��<�T.B�QGFbf3=�JnzF��D�KE�.��9����˘
L�'�rS�o��)Zp��h����9�J��{xn$� �O�e����y!KM	��t�d���ȼA/��̽���/��0�"G>y�f._�j�>=����n���^q!x��Kі�=W�51��xR�*W�������P�L.��Pd�G�oN.�J��5���E[����=U ��ރ��+Z���ٺt�GF{��
mXlxVHYEB    fa00    10c0�B�D\w���h�
rrZ��``��\������Q1�����<��R^qs���U�(�v�9�1o���d�}����	�����l�蛯^�C��,������B�_�_�q2�)�ݯX0C��0L�$G�R1����oc�`���+T�[�e^pV�l��곴�O�-ݺX9���a�O�M��u�R��ھ3�(PU���Heu[	q��W�<a�4��ѺXa���+��B'^B���㛶i���i(��͚��j���:ӞwUPd�������7N!��k�L�c5�������\w'U��Q��Y�e*$��!�b�`KVM���&��q�1����aYK2^0���1���x����z��:)>�1��H��t��q���i�tK!�K�6D��O1`�D��>�0k�/´����l��&�c����:��]�f�^ȗ0Uv�ᮈ��4D��C���saE��#��O�A����6�\�aZ�]xZw��,R����_α�X�M���_[h����jn����;��t�"���u�Fe�Q/h��G��w幈S���vǻ�� $(�n��r��ఔ:����Ln�dXD&f�%���0����fk��gV�o�v�FQ����K���� u7�2OI0\����B1Nϙ��6#�����n�C��=��c��+l\̃q8�Xe����V����E��h~:������,Xк���<�BƲ����@�	�CS�5;Pؽ����8�c��)Z��:�|�?�5���pi�:[�U�F��<~��W/�]�
@	VO��gJv���{�Zr��]F��~8�������r�x��/�.M�����+�Ge��I��R[Ƹ�'~\�&q������j�yO�t:H�`XE�����G~�	:2�_�?�D\6���	D�5�z�̥�Z�UKzς�V��mI�#��Q�6��D� �`�'[��$�D0^���׈��*�Cb�������a�W���g��V<�{����ב���Ŧ�v�z�1�e�/� �����5�x��Y�Sq����Kɛ]���I����D�\�WL��� �k�	큧�hC�5�\dq����z|zf<�^b�����j����U�{}@L�ϙ���i�-�IR�,5Rn�[�o_	��J��=����T�Θ˂{ޫg>�Ьlr!r�I�9�+78f/���/z@�z�#��#H����N/�nYac؁�d�7�M4���2��n�s��R�M-FJ+���������\�h�ϖҝS�/��똄�~�SiH����i.!0}�+�)'��Xʷ)�QT�?#��2�!�>��#K�(�x�N/:>N(X��r��h�y�� ?��>j"Q����2��*+���;��<�}=y���3~�<9hYn�_�!Әiy��8'��_~����2�k��.M���u����p�V��ķZ���{�i��
�\���&�UM�/���ZV�'�~�PVB{mq�ᶟH�@ޘ�#>T���s��O�3]Z1�JC�2,�|,mS ��s�j�\�D!~�B<+Õ`�k` 6w���%*i?KX
~�ܣ6꫑��|I�zuK3k���>�lN��wq�)��=�h���5U�
*�q�fE��@D�����3Z���W� �L��A��g*�wf�AV�Lh�۷7H-�#w�Ѹ��\�8 �'o��
��,Q�CXA������%������rVaD4Z/��{ɿ���o���駱���G�5�0Y��>i��^�����r��.��GGMϯ;/����~M�?�y�d�_��q�(���,{׮�qꅗ"��"�#��q���3l��������v�T���})�|�&��?$~�-O��tQ� ����±?op��p�M��I\�!C^��K�b,�k#- dI	�<�9
}tZ⢯1��#���o#�~n3�����n�p��;��i�J�
��1��A�C�>.� ��j���O^�p�Z�`��Gp��#���H�������H@��G��Yo�`V$EEB�&j$�w�R��r^	����1H߅��b��J�7�5V�I�7��q�js���!�	}E��/R��<�9��d����T�-�e|8!�����
HKET��lK�<�=*8�2(�U�Il�������9/O ���QFi-�m�	����e6����B'�Y��������e�6�h��M�3�d]�#�B8��J��gu@���SJ�̻nƕt��+�|j�V�{�������Imxb"|���NR6�_��{L�����;[}��"`%s1��?x���V	QIM�Ś��zX�NO��{������2(�e�"�GZ~�tWzQ�J��amjY��i�B6B��N���k�e�O?oߒf=�~Dk�G��ƠIp.���W�;������E���&���d��0��}S�	X�P)�&�w��AM(���[���������g5��^jC	*�Ѓit�[�9�m/�����1�	^*۱�A�t�;�K�����e�:Wj��K �A ��>�A�g'%~��f�*,�x8�0�?2�⛮��S����)�v�����&5\o��ҥ�D�5YN�AM0!���׌���tPD��+f?���`Ք�CЖ���ke���@���1P�"q�_Y��,���ޘ�tϲ��)�x��4=K*^n�� H��p���e����| {��T��S�}z�bNX��\����f���9$M�]h�j�!a��ԉ5`��W\2��~���٧�ﳺۘ ��a�M�����U�yY�C"����k�k�
$LP�F��X��v�k������ШӧX0qa����{� Î��{�����i(��"J���~�X�fHኢ�Hq��j�a�:~2��n�ts����_Z�"�8B4JɣEϭ���m.i#J��h�Pp֔��b�,��i�^\��n���~��W��k�Jl^�8%kO���3�	���@IЂ2M�SE*c�,���ʭ	��hLi�9��ö2�
�6�?�$@��d�3�	�o�O�m�n4.�!����7��Cf~����C� .�%2e`�)�F҃F����ʐ�4H�ӏX�˧�;������f9� 9��}$	y�4ZĘ������#����1��Ȼe��"������B��A����Gvr�I��̀�Q�����vC���Ȏu-�녇V�g�D�!g���B@J��N�R�����������Ħ�2�������g���efx㉶��+��)���V�70�s�B��H��Q�/��%�*���Tѽ����u�/��GI���Z�U��:����Dor �]M++0�}+�u�n�#]���n%���S�0^������b~�/c�_v���5���c��t��e��ΛX�H�/�����E��&�n�QK�%B�D��v+r�Ҧ��9��<N�ʨ�9�a:Hl�߇�Ic������(!��� ��b�(2R�4V޲��Q��ޝf4�v�Sn ��RM�G����Ρ�M��qh��[���4D:Ë��َ��Y3/w�2D�
Wi�jz5VT.�M[eb~�������RL2�N�m;1X��g�l�5�Gch�lH�T��4��NX�����'HrY|���C�6��)�"�Ǉ��~(��M�V7���{�iŸ���x��kB5��YC�]eד~7K����k#bv�h*�!���ed=�|g�I��{�[��f�Q�-[ꢨWY���˯����t=��C��?�#���XWV$).l��.��q�k[y����#�\�6b�j���eLNub׌�eW0</z��2�8[v׹�L +%>?`��{	m�Ԯ������*X^l4@���>��H�CJ�,ܭ��P�Ed�h3�;ͣ� �����l��QI�1�l�b�ߝ�?m��-����=W�X�,&-�څƿ-NI�I0��Tw޹$�m���7�w>�V�ƹ�\CP&|�[�^��"}j���A�s����K ��%�A��sM�:��^��Y5>�6�"UJ�fr�ۊ��W��c�E&,֑��M�Թ�
��%�
샲B��2lovAq���A��k�e����� �`��۟)�
�>p�|bG��?�@.��[�N��ִpP�~���_yx/4����!u��eă+: _����/ �Kއj�f����!4�ta���wSЎ�N�\�(��#V9x)vz�6ɥ9	1��ov&�O�Ǹd៲�e?h��Lÿ/��XlxVHYEB    fa00    1140�3wvN��/_P�=����&o��d�u9IX���6@Z���]'|�]�^��#�9�|�Q�0K���^F>��n���'�LI�ѕ��)V��.qJ���?�؝���/+~Z��t!��F�����N��AU�~!�����qb
������ ��k���=7⥑�2��
 ��8���-غb�h��@�G�c������s~�v.?��z����s>�\H�E�&�RNb��9K�վ4�g*�`�̯�P���8 �/!I�,�c�Ww�TΝ�,x�'���R�׹u΅�����ؽ �L�����nJ��`P��6
-�N;��ztb&m8�[��6o��"bD-Aë�ٽ�; I�r�o ��
"3�<":�LaTឲ���ـ�x�b1~Emw-�L��%����y%ٞ�䁆!x��lڶA9��z�i$[��Hz֜)1�����{;r��V9@�R"odo4�Â���Et���J��q�Z�t��!��$J`��L �ޏ�Nx/x$U7d!�"DZ������A	�U�c%"�n"�l��D>oK��+�X�������I�fn��\�R��SmqP8�����,����q�K��Y��a4*H�NP��|���}�A~!eK��A��i����Z]�ӠÎ�e���Ix� E���:���i������-�K&�I<�08��ۻ<���"8M�p�|� �M98�V^&�@���_�I}��L	�T-Sm�9l��S��0��YO���߃�b�>��w�j�H �J[b�	��Ð��nД&�R���^3��%��r]�Y�-`vrR�T���!1�����)#���v�T���G���ЗTH�fdY��$E�"6W�'��6�j{��P$�������p��}�����6Q�*�{�D>�T=�YW'Dq˙JZ�d�߽,֞P���r��~
p�2���|�����.f��]e�z��Z��~X����@���ʉN�1��R�P�<βڝe6�g��L��]��#r���l��ÓAr��#{�$�I��a������!����ѹ�üf�=t9���W����7�?��Ѻ���v%+�B�p���ۿ����"����V\E�v^���YA�xdx2T�YO4��祾���UߟkkYB.l@60��� ��{�h(����TEG���*}����c�=��R�l?n�����ް�1ӐM~!�sA��Tˍ��]C(޽����d�+���ut�V@z�x�ɔ:��w�����R�i�Z���b�F���v�R/(���!.\��`F�?/f_�b�,��0�.�.�:��1u�V'�KgFB�$���,�=�%;��G$گ�����C��q��]�k'����I��|���7"[�䇞�z�\wH�H�7�t!����Ya����<���Rs�!`�b]�\a����q=Y�w"~:��D��޶^�圪�`�ȭN!w�Ў Dnf��yrJ��ʩ�EdJ�]�uMJ~5`���>�����Leiub��Qk�aε^fL*�-O���p|)�a.jׄ�KcS�I�ne4{-K�s�t[If����!Di��;�^fYg�{��ٗSJ�$�N�Wo9I�x���D�в/R�;��܉����nC��}�x�y�o�7�zH�D70��c�X:�#�d_�/м9u�!��U�^��B���O�`�~��aZr�0|�(K ��_ ������u7�zM��]n1�L^1��e�nv>��\G,y<�(1�=<�790��x�V@�-�nׄd[wv`������Vd�
KP#d��!P�o%���K��`�=��"¨^�)b"q�G0_�\2>Dc!���2�1��[� %�և���y�ʥ�2^U͓��(���ݩG�ۗ�r�Z̆X�Y2zЇ5]_�K���߯����	�3�e"!��:�O�2E�0"a��-�|�y��x޽��;�^#���3�?F4<J.\��#R��:H���­���FRO��r�b���ɖ�����~�I~�&V44�y�]�{�T ���2|��hw���J��L�9�i�%UfS���h�G�?5b3�� �rQ�z�#-}���U?�b�fn�99t5�����g���>-��w%ȑ�������9�����x����B'�.kjb�`�:�����o�c~���X�u�MU�q�ؔ^���t��]�R��f6��q1�]�
��x�B����}�1���K�W2X6	�.T��/_Q9(c�ى�pE�Ϣʢ�AC�cPG�����]���&��;p!�����/R2_m��s����3v����K���	'��݃j 4�@���f6h�g�S�D
���	R�+���"�xz1r�0�C�I�����O���/��CZmoE����2in#Px]9���XF|���*>P�\F��{104���t�s~�����E��MrO � �(��*l�n�e���ƊyHy-�^�	z�r��ݻ�gP+g|��3{ڼ��p�R&@=p�dR*���^8��Js��5#d\T��	�Ta�t�wD;�y�q�&В����h�J��G��&R��K��L�0fQ��U^i���V��|'�^k�3n�5���1ı�[>M�S;T��Az�K�}>�����跕+��@�ž�����O�t}��U;�I�� �3+�N(�tWf��݉��6��k��T��&������T�����ʿvZ4�z.���q��΁���	���p[i���(^m���ʢ��� �3����%�_����ki_xՖ��8����� ��V#�����������*�U
 qT��AC���YXK#.��^�s����&dx�[A�m������1h�ل3b����ȖewN��L��������> F�q�X�⯠a��,�)��u2���c��״< �N��e�>�0��3���$������>I�[�g�κ�L���>��˄U|�0<|#2�����������M�NÌذ���
��$%_�>�p�4�?�?�9��dO��v]���uU	�ξ����Q����M��cfE�p��x�_`��d���s���_4GF~��7�l:�*�R�0{�����	�G<x{��:L_L4�F/�O࿈.�3��Wh��~�K�%��^����vh���b�q��Ja�|�#���ᔷ���b�u,z�GP���!>��&��(���7f�7>�ZJ���{>f�����k�ּ��#����eM�	��u&&�`���~󭵆ty�����8��u1�`�&h�RYj�k�K^�9<P9-=b�g���z�)��S��V, ��y촯��f�,����lZ����T��,�,Ϲ�nBC|���N$��8����"���qz��-�orڟa��t���s�o��3O����!�$f&?��%��N��S��z�g�W�@���@;�['>@Us�eg����s�sk�ui�*�^@�moK�b|{7�p��"
� Y�N'�{��7=�d���GW�a���B��:}�6�4v��t��h�?��I\�{R&X8���;�}fX�^��6�V�uwX�c.�0 �(�cS����}0M�UL�k�!"�����fM��0/�_4�A�OM8�z�W`�-[ta�FClCCC��<�#L��"G(ߊb��������(x��
��G$���n�CA2�l���a�J��@�>7	񆚡�?m�
�* R�"%��2�W�c��1A���J�Ԩ�#TrA�r���L=�戸�~�f�(�K�ؘ�\�u/7w)����K���W%%�WY�i{Ŭ����������Bޝ��\��Pg1�� ��F��/�v'y�!6�l���С�#�6@@���A�r����{E=�D6̣HO�7�CިԤ[6�h�W���&�X���`8�#��J�xc�M-wRf0��v�����B�Xaa�<VT!f�T3MD�֮��� �?\ ��&Q 1*b��E�5@��̟+�4��vI���i1��τ��@�#�I@�"���%#�1�ʰ�$7�%�����3�(�٩���hSy��5r��BS��1��/���N䄕�'�]�R�I�+��q�I �[uI���F���!�5��/Xf�d��[5M��Tu?4�ܙ�}gƻ��,fe9䲯P�}}qY�������r6��Ԅ�-w(�n�7�nS,"5f�xi���]��U�_E����p&�){k�6�-�+'u��:$��£R�,��H7�ۿ���=�� �E�4�����"�O�&)d������'5n��)}P�Gt�U�����1�O�ρ���efZB�z�$���i6D�K }K�zOA�]X�*�L؀�u�(rXlxVHYEB    fa00    12e0t�;����Ⱦ��萃S\@��*l���i���{�L0��-竇�B<5N��!�fU��60;˒~��|:�~?�6�� y�����/�r����:ȭ��y�1W��.��<Z�u��W]�;����þl�k�zm'�9�:��9���Y�`����8�S����^��4�gq&j��?��>�\�X(��S��)o�m����f�Wj�&�j55И���3��F�?�E���}��3;�az�5�M�G�p�t��]g�z����[בDo���!�i�t�_s�����;N��|\u��5���)z�Rocq���-�9��BCV���2���7�U�|݋�&�FMx��f��h��0f��KY(�F�^I�`)�R��T���C��or����_W-EG�8b�d�	�h��CcU�0�{�#I����������N;��t@4���
�8���d8��O%�D:�x�{6a�LNd�۽_�v��� �HU���'U�r�Qg����1�F:U1-���m+W�_���ZLV�qL�[�«��ڪ�:�!�p���Wk����4�W��[�5�����\��Uh#���G{̙�A�~.���Ė�C�ޕW�sf#��.�����f�����̘�ǕВ�M_v�Y`�������|ȍ8��穧���3Y]�����	s����٤�t\�	j|��4���L��	������7�!\�l�R.���Q����Q��}���Ʃ�6�RK�P7��'��A�^�|�4�	5��?!�@��6��	+�(��`̈�d��$L��*'��ؼ��y��6$�p���fr��{P�$���O�^X����*p�E����Jo��A�4�.�L�������8#��;Fh�B4�2��,b$:���`�s����A���ϽJ���x�ld�'ڎ�Zj�����G�@�Ȼv�c�,���5�٥���/��8]g,�v�~'� �f��)�0���a��b/jבBH��Y`՜ 3����ɤq�Nr�C��ٜ�d6^�7K	�K�o-�	C܏�q��������t@A{U?�k��Y��?n����f��~��z�eW^�}�hn;���������K����I
�آ��$�vr���u�(XL������z�pvqgH��%y�=������(���v�P�l��>S|�@Y��$�C�u�.�u(���WQ�1�ׄ唋7�˕��6=�tㄊ�Gu%t�&��(l�FN?t�5�jT��9��&X�S��:n��J���S$v@wv��:���)}/#�­����$K�'sl�u����j�|I_q���_e�6�s��$���N�0:��a'�����֏8�&�#�㋫��>�=c�>��z�\P���G�xYTYF�����Kd���D�M��Scfe?A*N�����j�RG��DƁ��G$	�u�mD�yC��Pk=��c]fU�F�\M�c �`p�0��*�%va��~&P�Q��9,��]����Z��&�����]�}��`��k�cV`-4q�!`���ԥx;��V��VH���1�}t��Ż�&X��6���)0+��Om`�*o} ����܆%�����/��֛�+%4�����X��U��H��t鏋5�r�P5i^aݍ�k��Ѹ*$wz|3�FJ�������9a�3H�U�%j'�Fi�88�R6����$����߱%��ǾY�4m8�g���C�l`� �8^�ל�<oXu�n�~iY��^dZ^l�4��_h�@���ݕ&U���%�i.+�K�E{s��gK3�X<;�S86".-('��?�=[�l$(h���~'F4�fQpq�f�08�Ҭ��r���K�/i��&�T�E8�>����U�~��~�UFeP���"�W�ٸ��S}Y��[��!V�ſ��|�yp�D ��S퀥��%�iw��d�`E����^�2���w��[m�x����}+�/h��i|��_κ,�0|�fi��yxR/�����âQ#>G�r���bQD|P�t�b�u�4��������])W!B��;�ް����}����S]z0cC5j�T�����&R�i3�	[]=Yҫ�\����+>8r�! �4�8Q�;�xc�`Q�ï��y���9D�K��@��2��<՚��<"�d|�J"?^c��(|��D��3L����}��o�`L��~��'&ͻ�d�U��z���2D��_��$^l�ě���C�q��ڢ�ո�FUB�D���:tH�;z9Y��.�^�\��0�}�W�*�+�o۠"Fj|wI���2M������PD׵Ao�`ޫp�$�7ة���G$A��@ ��#:`�$
��?�zg�[�0PV&�+�UY��\��/��B���G�-�f �c$,yD-����g|>�u�;ەF��t���sI5��a5���������EC�	�k�$��)�GОN�V��R}�ِ�V��B'yr(?�f�M�	�Vd���B��0������ �����3|�����S0R����Qy��� �H{�{�^*�q7�j�]�eT�^�q�l�����s!B8#���7*��)��;P��Kh�����<.{���Ѹ(!~�|���uF�-)��)���fK���ù���p+3�ɬ�k?Tc�O�*�'�|ƛ��{��d�����"��ڏsv�-����Ѝ+�%�)`wPO?#&P\h���D֤����~r�)�2�i���/�1��9�֯��T4^�P;sB��	BCkT��(���'3!.�/�W�RE1�| �h������]�'k�R$��qع�'KD)��/�K��1��v[+;
ߠf���z��XE�4��j�z�s��ىo��z㸡�ڤ��<7y�"�%`�d0���8�*|)��f+�,m�RGY���,8qv��a#���jZ�]����p6��G:�d��~��w�:��
xWx�[RȮ�����b���vz�MD�4���Mar��ag;���^e_��NEt�F3����Y�?;>��FC�ؾ�u�k�z*�Zn���n������ī�?��^�P�6
0��DڸX�p�R!�c�t�{�W���C�2�l{L6��mf�/I������,x|2��!H���
sK<�7�E��,�cO�+6Xi�=��-@q�����%χX��<��(�B������U���|���.w��<�94ʥ<��& !
�����F���U��J�v���\���Cas�7��p�F��m�6�����f�%���!Kr��H�e=���K�a��Op��ș���x���-�qOb�}Għֺ
���F����W���Y,Kh��0Y;#�j/0A��%'6
$�x^*�r�-��Xk�bq���{��^��f��o�
N��+���ש@�s��c�x/�f+�[~�f�'�'�v�!�E���ܫ�1�  ���0�	�o]��]�(T��+m�
(@h��{��.�����\�2~O�r�69��)���$��J���߀b��ط�W�К��	�zGk�����&պW��,1w�.	P� �璙\�wRb1���X��7\^���=��1�K�RR�a�S���Ŋ��$K�@�k&o��~�6�SC��|]��S]C��|[s�}Õa?�ǔ/�U	z�$��_'g��о�f[��}*.�_0���zr��[�R�M���NR�7C9G�U|���N���a�UxM<&�*ܑ�����Ŋ�x�Å�( mǸ;�F�Y��;`#�D����HɗM(F�F5��2�����9��u��4xoO0}�8�
�Y�4�/������l��q_.$ ��mHI���y�^��l�-q�P����뒱Vs����~�٪�I�O5�Ck����T�<�S��4>��<�g��ن|vO9s��i�ɻ�\3z"�]�ɔ";}�*%�2�0Q<�yn3������5�I�ޝ�>[���; ��������P��▶��Ӱr�t)�&=�����k�����
�j$�`�%ix�m�D��5��z���'��.AO	�ա�����B���%�#L\��m����9�^nn���ΰ�ę}�� ���m�ԏ���"�a�{� $��J݀�@���e\�$&���W�8��{UY��顊�l�Yw�%Ֆ��X"z�i�^ �5�9��D��+lٴwi{��F퓐_�,Y����g�� a?CC�?H�ǲn#�w�0���ަ��{!_������T�w�j$���Kyo'FjP���VY��!��4=��ZN������w�$G���4��݆{���"��#m�V4�ϫ�e��F�ShImn����������a��&�̨��-]�C���qX�F�f�l��
}C�Y����g�
�qo�nb"�fB���ߗA�v�T�=�l�"&,��|Y����R��0Vg<5Y��)�\R�[���:�j�'���jM�d��YAr
"')���o{����e(�,-$���3�r
3⠱ƼQ�`d���ܕ����T���]zi�J�u뽕JPhո�U�h�IkE�6$���x����9X��W�q^�V*zd�C<��TX��H�	��/�j�����L���+̞yZ?�J2�u޳��<��8����>Ǝ�}�\���]�����:�- �R2�RG֎�3#%��&��X�c&�Md��<�i�y�`��l-eב���G�1V�_*��a@AS��_2A�l�6#�O��p��ܯ8r���z��@1�u���~[�]����XlxVHYEB    fa00     f50��nf3�4]!�XI����Af��|W�𹛦A�D�bڙF��}��F7!W�1mk �ċ<5�u4яR�`b��
ݲD�҈8@����7�\Ջ���'����^J����J��"�ZBR�κ=;��v.;�sW�S%A���⃀��`�8$�D�}�H$�(W�)�Ӊ�#Ez�P��I{5��%&�%K�ſv,��H\rɝ���ެX�S,���o�d���ҽ�b�p ~u�)�/��^� �W��＂�?#���Cv��_��*���BH��+�gj�|N����N᪶��j�?�5�L�=:K�M�NF�5�?����e��E���e᝝�gzP)L%��9;��B�U?d�3/�����P�ֲ��|��|��ţ� m>��LA��<�oZB�Ë}�>0H� �n��`am~D��,jG(��T����rdc�ad��ǔ���5gJ~��f���Y�����it���Է��l0gε���%Ƨ��_��Ip#�,�ܠ7���3`ʌ$an)�ܗ]�R���ј�O��'�'�^M̸@.�>Mz�������ĞNm�d�r���6{��][l�c �ؒ��1�fm���D]-|�x��pN'��'�o����&D�H��1�څ�� ��pW%4�����E��颙JW�Ap��D�ٟ��x�w׸�h�v�o>p*���=y�,�3	��=jT�Soj3�2lq&)R���������� �pZ+�ʟ��+�1|�{�kݫ&�cO	��ĲO� �й�!�6w�(���@z7�"s'�~�8�!��a���7��?t���(���9��B]�r�J�gq��Ů�ʗ��[��:Z�y�ȦL��$k� :�WZ��Q|c�,�L���U�o�U<#�7�jZ��?��)g@g�E@)*�J0
��wb�:��ϞB\>���4o̺�:�6Ȩ�(ŧ �m�b��V�9��_�}D��8��l��\�W-8��>.�ҝ~�;.�;�z���L7��=Y<=bs+gT�
;=��d x��̂|=�O��������0�p�%2�t�=v���(>'�_f�?��P3o*24Z��N5�G����آb�f�3�#7�,q�?ա��3��\�V�T7z[����"��@&��]����Y�8犄k�R��O��ڏ�D"軼L5��ع?�o:<�	���è�˲g/�߀�X�q���|���-�')�|�ьo��Q&��η����ю��6R'g�7(�X!h�59�5'
j��s�C���!6�	CIŁ"���+�R5�V��s�V���d�[mM���m�b�V�����A��Оz�Qss��*ށ[(����xU:�WH]}kg���*^q��8a%䜷���KK�2G��b4�z��>���p���/�d��0O��q��`�蜠�m�4���fn<�^*`������(��4�̉�x�������1�p���kt
��(p'��]�nIC������WU����<�=J���%�=	+���$�.?�d�ƌ�������#�{Q ���<��	��Ӻ]����1��Qg+��a9|i�`����fjv�,X ��6���<B*iL�$�7e�k�	��Ԗ�Y��9ݵ7Oک��\w�F;��*7�D�!J�-�M��Z(L�ܺ�@��v���R�eI��U�xk�I�B!�m�#��7��ړ��d����Q�U���l=/�1�af ����t�� 4 �IHW6��M��T�7�zu���e�zi˙H�JfQ��}a�xF�6W�Ћ��m1Mi��8�Nni��b_�Y.���P�q���,�"�N��ɥ6�[��NM���_��L�d�
�Do�{4��嫃�Y	c�!�{[�7\9a���}�n��8�/du��y@qOKO&5V�q�b�g�#��Js�U6�"���g�$⚇<������{0y�	^�z쏧�+�X����y����H�`S�P$4fl�nk,?���n@�eQOV& ���n۽�L�lv��� ��A_;����N�n��9l2m�\ޙp���*���:�s�2�l�T̻dkw/O\���ﴇ#CZ&n�f���#5�З��#��͡��L����{�,O��Z�3�Ao��>�L�V��^Og���&7����(�#����v�ŮҺK Ӭr�_K����	��P�Rdy"��s;��\vG�i.��%+�Nn�����#�ã�i�t���%��g��q�j�n2�+���@[ggEM�jB�<����+��t�d�0Hϱ>�H�v�~�T\N�o�ry����v��6��M�ϳ��6�
Ze�������n�#wgfUt�)�#�7g)kE��or�+(�/�(e΀xJ���ƪ�
CH:VL7�4�o���  ��h��*�#R�*%+KD8/��:w�z�y�(�Q|G\o��>q�㧆P�U�m�F�-����w}.�䎭�V���8K>����7;��{�U���2!�,jr;j �s�����
�X��](dGyh�¦�q�L3�v�:$�>1 Z��w�.uC|F�\'U���[�R���g����@����X�I�+����M����.%����g��m6k�_���
�3�:���D���f���!�׵�d �n��8�$��9�~/��tK��m6�`.k}yf�n��.���lI�)��cHqP=�'�����B+72��x�kz\,j�ڱ���_��k�$9���1i�[�w��m�7�1�ٴ���0�_ ��W |�;B�QM��y����q-2K �E��!�M=OZV#���5E[��]j��bb�#o���{���$��Ns�Z���F���:�Jv�⋇C�4vz#C����,��@�|h�x`���>:��)?�#"�K`s�櫣H�m���q���F��x�����:0_��������e�r�S��7�Z��gz�W�]7����7����w�q��Z(Ύ|%k�el�5Qh��X4u��g�qU�h��K���@(���{y	�?����][�?�*܀�����̾��f2o5�ɼ�7�CrD%1�&o���`�2+��/<Hv��� �s*s�Wj3�q�`�l���֟��� ��T��!5��v���]�zY���flU��5�ΦL��dVt/�ߎ�>�^u*�d<!5d7	i�aǣ���?8�B��-�^bQ��������0៍_��50�&\�B�Ɍ�g��x�v�=�u'.!��xH�ݓ�R]{Y��i�c���lR��3"�>/dn��RU�fM�VF\\��b|���Ҥ&`�u�y
o1�����,x��Kt�2�v/MEy
�F5]eT���ۅ���e��F��yX�����~�(c���n�[���F���Ӫ�&�Ķ.y�ݗz0�)��;�P+0#�01�p�	w:L����+P&Aŀ��\�x?�f0�:�k����޴lD)�̶%���Xe��g��U"㷳:?�������d�V�/ ��kzf��!>�_+�sV��^n��(��3�#�D��䫉4c-�x��I���U�(�#�t��K?-�[�ې�I�a�k�Jd�GǏ� "ڶd�N���_>b��x���vP� �=�v��ة^B���,.a!�:-)�5ɱ2�7߫��ѣ��x�Q,ve��3G%F�L��M�����6B2)<�#��x��:	ok�qfH�=:����0�t�R�VO�>�&o���p�5���O`�LI�X�o<H��_�W����iW��6}�h�f�<_�1�bl丰� �����tTl4�P	Ǹ�낑$N�C���G�O}����A1���u�04..{�*��������O'��Z�3XlxVHYEB    7273     560��Т����h�>f�ݥ��D\�d8�ZW,��?����P&L|sl�Ǘ��Vnf!�ٽޔZO�g��F�q"��p�!�J�!��2J��>1��w��l�7X�PP H���X��{�?^1e)�5c:��sx2P��i��K��C�ZX��y���oN`���\/iZkp׿,�G��E�"�v^*�lpp�x5��&�jɼsp��E��I>�%�����Q��@[dn��>����De�v��q�x}ʐ�n$$�"�'�ˁ��!|z�܍��z���b�Q#��j"�f����d����5��̷��W.|��b��Cz�!�%��d� Xx�#w.ڃ'�n�`�Ǘ��=2VTe��b��=9n۴l���w�dM�A�3�)�6ko�݆,�^OW���#���"~Ut�:F!�w�p�$�&���Á�J�/ ����a��Et=��l~�Zs���7|��曾��}M�؏��
���0T�h���Y���+���&���&�e�
٣Z[Hq%��|ʰQ��G04aq��1ҎC�gU`������
9���`B��Ü��;M�8^F���8�h�a	u���G-���?��u�d��m�w�ĕ�؂�n B.V|���#G�tJ�\��gZ���� x�ި�.^���M�Z�@
)����@���X���������YE�����#��ʄF_�K!{[K����((���,�/���E�-,[MB gѿ)�*}h\��N�?����pgD�$���'�ET�C2M4� Iϻ1�}p�z\��83��nӋ�N�dW�;[3"o^�*)�Ș����7�'�$Uﻂ��\�<�j.^�O�	��+���F~B��|�쓾06J��;���l�/�ܙx��;�	4;����|ۆ�V�����S����S�������[ͣu '�0�x��)?�b�P��!���5g�;�)�B�x���	j��&�GLx�ak$v�+�����LI�<�YF��Z���K��F�;�j Y�%}�O`�ٺ�ȾP���E�Y��	�W�L���o���l.�GH���*���r��P`�拤p5I^�Ky-�-0��9����*�1�`��^���
�Nn��\�<x�qT~lT�Zs��%��W��
������nG�����r"��R!��a�'Q;3��cٟ�֢jz����4��ZS[ԓ1�i��*���������4�x��%r�~�ٚ߫6v�n�05P=��R|LR�R/�����]�6�����i��!h��i��_fQ��r���B׏�>��c�<��k+������A�8؟z�N�=|`�WQ[��R�Ѿz�_d鵯o�9v��3f,�m