XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��1�?���L �f�
��y���7G1�~��D;��i*�%zC-��~X/}�>5��p�X�/�+��8�����7 ����摲^�x�5�
8�/�:ʾcz��X���|!���OA��*w�Ncؙ�,�Ri7��'Cp�+����5V#T�Y0��+,~�v�^,�5������-/��������H���{�7��~rj;0���@l�N� ��+���W~��V���@��v!�hYQ�טCj���q��D�Ï�$���@����	39X/�
���$��ʲ07�z�ŉ	����YG�L�#`-�g����\�&��G��i��eV���Ρ�d/��N0�dO��M�n� ���P>񤤳v�Ƥ�2L��"X��w
J��jSh����&T7��H���߷�Nw�+ʼP��Gy���K�+�JCew�,�Q����Kz��1���C�k�i����
 Kiֻ�v�r���WT�ͪ�["��6�v BK������#�wq�a	)�¯(R���Ȱzgq�d��0������dԚSf���	M�r-%�P*įP��+���K>wh'�y��$H�s��M��+0��0���E�b��0�����ej�٧~�� �b�!��#����8>L����������|PO��X����ò%��\w�?���b˷lS2?V9����7���\0�$.x�x��%�R�4r��� ��9��@�g"䔤0���~"��(�k�/����	N����nh��8�f�L��XlxVHYEB    838b    1770�0��MY��L?t.�e���/eܝ�~�X[�2��.�տM3.��P��\����[[��(�Y>���N,�r����Uc���#9�k7HOc�lYsw2CV�3�TI}ϡS�4�3��Y�-&ݐΜ�=� (�H�	ڕe-���gN�x 濛���Kk��Ƿ���΂K%m��=�7���o�A���,R�\E���}���0�T�5EV��Q�q�q�$Q ��y��W`�զU��~̳��9i C�5+U����Ijk�-����[rܹ���ɰ`����?@�uY�b�($�O7N�>���g;s�ͻ�N�K���\X|��!^�«���Д�|��}����{�� ^�5e�x�鼋�8��Z����,G'�+�/��$�{6���E���y���,)�����',��h�)Shg��6 :y�V��8��%�)R�fe3Ut.�w��(N�0h�_�n?�[:��%�e�F.��
G�hI��2���5�_��D,"<D�v|�A�\AN��W/SY�(��+��1
�|j�s�G�s�����Ȕ�S�\�k�ݮg�%��$˝���~2EC�HȔ�u�@��Z��K(�^��S�x�Q%?N�Y�e�G�B#�2ޱq�hϜ���^���um�#�T��"B��-� ��m4j��K�s� 	T�W��9fÚ}N7+���%�$ݤ$a+z=�� $�`9������6��_r�8�g*YE0r'���a��O�NG�L��5hS�`�r�ǃ��
��c�W�@\n���\v(�	K)�����c�<m��b�ա^�r8��/m�Ѡر���Q�����`t>��$7��k����޼�<2[�<w֝�n�������V!���Q�W��U�|�᧠%?9��6,\_7���up�V��Б����7K��d\�%Bjd�b��zZjt�e�*Fˊ������%����$<h� �ni&�0H6�/��1�i�������s,h�^Afp/�v�nͿ�L���5	\�O�3j�~�b�6þ(��C^���N��l�mh�-,e.�8�*��"�����m��0�\��	�	%W�ͣ��r K�SMi3��
�_,���j�O�S�%���`,M7��K��N�9_�>6��E�0��i��1�g��cs��A��Mp�5�LhwS�ߓH������O�.yj˔���M<���F�ޔ䖄�������	����O?r �³q=��wJ�r(��jA[�V�gf�/N�f����.;{���_�S '�@ ��}KvР�3<�tQ� �/�Y)\*0�?vsg6~���ƹq3����q$�~WB$�����g�����(�{t��`
�����H6����]A7>��«�V�x��M9�����F�+1,c��1/�֞(=�?���X���2Ek�� :oN�b��*3 "�i�e�|�M�x|�%B�����|��V���J.��R��,�L`�c�{'4�<�`����yH@>���**�C���(�Hu��$x����+���|��H�`�lu��B����Uz
N[V �U��j�.8����tj�N�E��~�ba5sU;H�����\�,]na�,�Þ_ �`�6��*�u�����_?�Oxw}{�"�Ox�ˎ|D�6��Hg��
>KS$��ƹ�t~~�}f��nv�t�QZ��l�?*�sVa'S�;8�q���瘼����g�>���j��b����;m*o���.{��(Nt744��Ջ*�ˊ�5�[�L�`�fK��;V��}�����P2�M^;�ZH:+o���d�x[V 1�����f��ʃ�i-vÊ��FZK�x;b�<�1Q�\��]zoV��ϳ�
pb�Gx��hF�pT,4�COT����Tja_=s���/gJc�!d�6=�V�M�gc����꭬`f�����g� E��^S���nqX�s�Z�@0�i
q�p�XA�^�
�.
����z�|֖��3�P��Y���'���G7[ˑ)]t�z�?T�2�FJ�
(��◩��Eq9UU��������(�n�d��~����L3��$fG-��5q�r��Fȝ?�
��3^2�1��,�tޱ,"�W�*��ʸ��>����tc����v���O6ύ�u�dDu
s��_Pϸe�J �a1v����,���4���~:���lxŐ���k1�|�ل��X��yC@�.�U%����GT]�|�{�����藞K$'������#�6z*uG�zb{5�rʦ��������:��Q��L#G�ʈ�̎c�'�W�ǣ�K��@���R[|İ�$2"�~R����Tڟ_��NM!e�lZd�Fu ��:���p}eV	�Yzs��ŋw���u�Glh��G��Z'�^"L���\�A�'w��X-Z�u#���_��	6G��,�`�t��a0�xϳ4���.�}��~yGy��`���M/&)�������N��6��u���� ���vy�d��'ۦh�<!��Ӣ��<f�|��O �Hc�Z z�S�󘸇�/8l����%�u�1j)8Q�kۻ:�}l�f�?���s��1|	�Q�m]p^���\HTI�t�}�Nz-��c���Rˢ4ɷ��L��R��0�F~!H]���a`�;���s����m��=G�mߛֆ�K5s?�Y�j�tF�V���88�\�j$��^�FSE�2+��M��X�!���t5�-W��RK��)�[K���hHQ��B9�����=��:؁�$�w�V ��Z�>�0�Θ��6��{f�����s�	�6����P:'M�c~K0JHm���Z����B,�!�I�����^!Ly*�I"�YC�b��;4���r+�g��-�b;Z-��ok�vd��8��Z$��m'�7��YWt�bv'��/�|F�&�?R�%�Ъ	��F$���?�94�1�e�F�U��Xe0��03nd�=Q?�fw�:��R�&D�K��HoD�n(��X�b�*���}%p���aW��|'v�FB�"�^�Pᵎs��v����Zsh�@�AU����d��&�� *���5������<
�|y���~��5u���[麆!t�e@�l�b�t½�O���N�gD�i5-a��KZ����O̉r���V�k�2�,��Ӧ(����S�"?��ym6��]��6��.�m`�gJ��!a���]w�`���e���t�`^��2�0�t���a�ǝ�����m��oD�p�(��v[�lp9	��A1_�(�2LQF
���ޢ߻AE��~��"��6�t&�Ȍ�>C���C��L�r[*1��,͜�T��4ͳ��&p�.vKᄠO��`�u���)3����i��q��#�\��
�E��6#\O�g_�����*�q�Pg_�sI�'�wqU4����z��٬�[��wg8�v�t]l6e���φM���dՓO\eg�ۋ-�D�.��VA��ɍ6�p��U�e��42�Զ������GIŎ)��<���<�B��{��\����!x���'�q)�4?��A%B%<]��ӛ�-ք�����+���Pl{'������Ft�PA���&s�����wf!�=H&����oi1dS�����4�����d����?����=��=�k ������ۥ�~�#%���P�)�@�t�G�RC�N��$�<��]z4#��q3�|3����7H2��b` �����֐�[�#C"���;s�iT(Lف��k��0S�1"�ϦA�·�D�9k������Hf"}۹��큃)[B�,2j�����db;��!+�=���03���4ݩ*o��Ee�0w�Z�Z�� >��R/��Lz0]]$-��/�l��k�[�ie|!�LD��h>Ǥ�n(�%D�&�9횦�8+L�R��"M�-z�3�^��8p�qcWq���:	VuM���}��	+�#�Z����	�~�`�| �r�~�N4�@�&��{�<���oak��e-�uʜ��E��,�c��wh��zH��ƍgn�[�r�%�&ZZ]^ל�V��R;Af�?8�L��-��v��2�\���㢒����]�J���f���V�p�f��:u,��S�x�d�nV�~N���[㧀\Y��(��mđ�i�"�U�L�L*�[sl��:��� ���|���@�'ۅ�@���
��,H����D=3G��S�W��z��d)�n���htIѰh�gp�W�$�A,��x��eQ� lY2��	�8�+<�/m���J;�u�(����ᬍ�٭"�t�Ž�3�ͻ�@ťm}��L�v��Gwz+�r+��Z(�@;;:N-�bcW���%� d�`siޛ����f?��	Eg�g��~�V��S�z����JCtF딄���ĝ��g>ZiG])7,v��yt�sI���5Xl4�8��'-��@*�*�F��$��͐�ICV������Q��ZW}���&<fB��<�qB��(��xD`I��������sP���VW(�P��'�%3�������lamY�.�V�gJ-K��
���p�����g�~��c�"��W�W�b4s4��XBCf����E�Jc��9��l�d�T��!�_�����	BGc_Z*!V'�o���4��̀|$oL鶮�k�'�-����zஇ�3wAD?�
^g~,����GyE%���=L_Z$��7�&!�"U�d2�S��R�P��k�28�0�~��ѫ���l��l��"?6��rd:�Kg٪��T��@��(پ��}�����k�y4#)�]�~叮�SM>]����,��)��OG����39Z�|:���,;PGI6�o�*�df7���bv7yb�I�]��>�"����S`�@�3p.VW��G<�������[��7�����8�@�u���(?�G��$(��`[�w�]�]�?����L����* ���-��op�,&!U�҆i�d����ԑ�[�fs0bB�	�$�
3�1��J��qj	h+[����6f��_��#��!=�R����S�uC'�B/b��o���2�q��bZ�r�6j��\�>u5�O���W\E� �ᢄ�r��ŷ�[��������`ɐJ�޿�i��w��.���u%S�?�K7��Y�n���f��2�����)lr��'�~b'��������\pv��l�c�Nk�N��m���E{�]����.`1܎�k7>EJ#��M4�`/�����nz|���m�]�Z��Z��s]E-�ƨ�Hж�1G������,��߇����R��~_�B'���5�3��zDP��L��2}�!��V>�n��%������ˇM|�qf0H'�+벦��x�������dq�cY�h�~!�|��p���M���K%�E�LlK���˂l��x��MR�y��C�}�3L2Y�溽~�<J���%_�L�7��d���!��D�v!X��>y����Oc�E�8bi��ˡ�D�ɚ�!����y;,�,x���ou�����K��1ĪJ�W�Ǽ�G��b�P��\�+"�~��"F0�㉁dܟ�Ӗ�]��=�1�3Y2r�ʻҶ|'��U�E�l����q�R.k{e�ǵ8)���U'R��0ڭ?�`��6#���`fD��a����{��٧�U��	bL����:�TZT��QX.�J��l���Ol!9 �Y��]�DvG �7
ne�'�FZ��j�<!j����z)&n��Y�Q��V�
�v��j;Z��{r3���������Op)�@#1�����C�^��W`��W?vi��IpH�w�X���:��9ڍ`��J��
��&�a)�h�c��g6���׺	�D�xR�φ�R�;9�5	�Z�Д��-�G�ϵ�a"b��GJ��l������d��O
=y��z����tP]���d"�b��rĔۺ[v�JK��C�a)