XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����E�$� ��Iq��{��Wftx��Y�@q��qQQ��P�t�X�9�W�7�p ���䨢���� /'�|���>��#)$��N\��<�߼��m��v[��("uץb٠ɬ�)@�zX� �������ش����8��5�A�>'�xgHU_�u�	��-�% ����M|ݢ�icb��CE�_e�!{u�Frk3��5Eʴ����&D� �茹s�>2��A�z�#�:�h�(��ME[���l��xK0�T�7=��N����B��;9��)ߌ��(x��ad	<۵D��@=6퀕��Z�'�d��c��=��t�)���-v����3�B�l�����GAхS�~��KI�s�|�w0���y���t�\4%Q9���l1��)�kl�-cTd��S Mti켂M�ֳ�8���W�A*���F�g�o�l���� �Ø���"�P���Q��R)�<�!����P�~ֻ�5��%��hKC�c@j�����A��W��FM����c���=\X���μ`�3f���]Tÿ���0�6��W��O�T��$:o��_G�����r��u��[LFf44��h�f&���n��r��
(jo�>N�}e�����)p=@�WBV���'��n�jO:����?]���q����Q����Eu��]~��u7IES�JQ3A�=�w䝾�<���6�<�e�^�/�{�C{��>��r�m�/'.�JC���u���&�S��Cld��<z ����XlxVHYEB    248e     9f0[Ea(O��o~cIu��`��a��=~�NZ�<�`)f��~�e���QW�Gf龴T�s�+�fb��GO�Z.���P!ͨ��.�D�`��`5�����A+�21�Ŝ��k3��F���{��F��T�h����}K�wf�4mIڦ��oV^V)�U��Rk��O���$_W�>�����h�?lr�ʀ�?���i��l��z}Wsa	l����v�N�u���A�F��]Tuѹ�dm�6�`��ml-����)LX%K�{�����u!��bVx6��w��vI �&���]�=K��q�6���pa��p��3J#t����1�kȻ�(ae�`~d8v�Mz�/���DG�K�$ ��BԄ@Dh������5mBUp��G�QF��u��[�T���`�U�A3��I
��D��y�G��_½zN�[	�$��Kz�ů.���b�kSp�N��L)��et<�	Vj��<��A�/U[�w��ɼ�re��4���ë���+>���
҃��̝� 5���Jy��1�0E Lfi��QQ��aC��k�#_kuzf�M�硺	Tﾗh�x-#�z�)	j�N��=<p�v�[�����AN���y�?�xq��}aC�Y�^
���!��#�&;Ӹ=$ @����zO3㵜��RP?�M;+訰�?��,��TcC�[�>ҿ1󢐍p��,��O�0�5�c�K�1�5�&�u]����;��O�?��C�K�l�]Qܷ����݆��Vh�C'�Ցݮ��ZY�2�y\�RI,jr���2@�A`��o��{ʂ���+��d�3آ��dF&��.��~��(4i�c�I��yh���|��$ݞ�D�"Eŝ��k6-�=B����Oĩ�R��p�E�7Y�j�O"\�A�,�˞F����|4�Ŏq�K��9qP�Р�w�-+��u���HS𘚎�:�,V�G�U�|�hN	�����;3@-f�us�M�<�%�$��nh��]O��M�K�0��|E+ovT�����x�3(���E�_�*%߾݋�z���I�7�
��t1O~|��EtM�t��V�ˉg�v��žYF>_���-o����y$n��I�s�%���D��j��$���� �0CB`:8ɉ����)�	�Q�������]���B��b�W�z)�Ɉ�uC�5iԠ�����F�w�Ǎnr4ک.ᗑ�G�T�ƴy�-�Z&A�5��	��Y�|A_gX7�yLR�x�6�4z�>xOkùy�W;#�7�v�W�)C�JL5j���f���Bs��uB{���4�]���5Q��[�c~駉�:A����L��	`=��Ȣ%���f�`P�A�%�E�~������Aύᠤ�?�,}��dA�{.�+Я�(y�\r���DQX��oK�5+6C/~�g�5�\�u�\�>C�H��GWB�������W�kʔ��Zn��[8[Zd��=�/3��f"�k����	����V��w�^G�FV�~^0�����ms���"p�"���?g�;���C�W�`�)����Y����b�N��d��,�;���4�3 k�E6Q���R���KǕ�֒�~$>��ͮ
5����Z �"�d�'�G��:�]l�>%s��0lz��c�`�fɠ��^`�;�Ԥᤏe�V�pCڋ�
פ:���7*G�`�'%ʁ@��;!Ţ�f�Hg�l�'yol���Jݛs��*�����3�C�$� �尵l�5��H1R���(h��4�Dy�=�{����'�#/6�Yc�qJ��U>{D���A�� ;=��A����͵avrH��<����qk@���w�T��f�9 l-��N�(�� �&��7 }�>-Ala����j�#��M9ć�7��z��Vc�N�x薍�SJǕ��2z�^��<m#dpYE�dʰ4�y��i� ˡd���4:W?rZɊ<�Fx���w��H��{m��|��xPEx�-O�=�i	0�rc���;�,
��	���x�`����VI�^�m|�w-N<���+�q��L_�I�D����m�x?�`T�A����/|��vg}~ҔKvZVk� q�<߀�����ο8=���h�������MR@0�~��m�R^�煵+`ew�T�y���$�S�\�i$���<_��
�J��-^tVܝt���	�p���"�'0v��|JE�έx�o����.f�����O���AD~��o��-���Y�(�{ruԙϴ�W�N�Z�k�ۏ�P��ŗ\�RQ
����p"��I�Q4s�R^qS��* B�Xp�R	D��a������DZ.�����>��LW�
ؓ�Ou�"���2У�cZ�����q%+���A�'�Q餚�@��TFJ�	�<2<Тg��!6�A��+���`E�f���2�$�r�J�]-)}���}��Y8UN)��g��H�=O�Mx��ػ��uڂs�Tp,5: ��@KN�CJ�9[*���gE�hv�h)?{&��ȿV���s�у���b�&e�����Ö6#&��pr