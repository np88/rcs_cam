XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����\'��Y�[����f,�c׽�Ųb�Z��!"8 	5�n��Y���Fwv�F��}J�S��s�#r�����I�m��m��{�u���wOR�9*
ĦT��xM1ߺ�᠅�=|�����a]�VY�A��QaŉvoѦt���
�`�E$_|�h�f]ib�s�2�fk��J�Uo�e��iLf�ij2���Y�姅��)K�;�mV�f�;ڡ;(���q�~ߥ�ɪZ�S9����ʿ�ALm��բ�h�z�ذ��`�֟�޹1T�����Vwa���ph��0Sd�	{5Ч���X��m{9���?�1����Ͼ�䝔o��g�J��5P�@��5�����ٙo��c�VU�WR����$��r��݁g�f�`�~�j����f��F`7T�R�x007MACA�(O�6+F|+�����/E���|�ـƑ���Ck<:f�+�W�-��e�i��Pl�Z�j2�d9LU�릏��bM�`�(e�*E��$Q���E�\��ʛ�Y9ّ����Yw�Y��Oq���% c��WȐ΂���%���3�M�\4Uark�VbG�R-T:�)���!BY���m 
��h�7O�^6']���ߝ�D���/ӝ��4���F���A׋ܢN��J��df�^��>�0��J������]��΍L��&=�����S������Ҳ�b��y��"m]���l��~��ѯb2��������e���v����9߀��W�E\��XlxVHYEB    1427     840�e��L+t?�9�������h���i]����8������qS&.�l0ћ�@~/ �esŲ$��jI����B�JuT���zͰ;mo>.���b�(wh�&��+��B(�	ه��Y��ؿR�׿�����\*be�]�in��& ������\}BI:̐� ��_��('�� �-���F��,�<^���:$�h_pE@_�����h �x�J�����偙�[4��/���s�� b��p�,���oYT�8
���!��=I�(��KŢQ$�D*�B�h|C�&8��T�di9-R�ܿ4�e��nI����Ռ��$j�@���P~N�ŉ��M=�
�Y��qOd�I%��{a�@<�D�n��ۦd�t3�/ʱr����N���م胇�K��Q.W���x����u�_]�X�ߗ�t��3�v����!ʤ� �EK����)����y@tz�uc��?��a���@�i��D�q'3�hm�,
�T8��֕�e|p��{�l�ZBw���6`�"Ҍ���4Q���}��AA�˩F]����ww�_Ԭ���N���q���)���%���OH!�A�v"O ������X��e�g�k<��}"~~l�i���!�Bo���x'�$�{��b�p�ra�uQ�g`U���w�e��f���w�f(3���ɻq;C��#��Y�N�����{��%�1�^��x����b��Й����~������}4a�6�?�����2�1�d����k�6IFI?a����O&w�Y��y�KK�8�����E҃[E*�G���q����x�یh:�a�x��e-=�/����>b"���v(W/�rX%E���Q3Ms��v�Ē��.�0x�P�~!�y:�? �D��FK~����Sɫ"(,S�$9���h�*W�h��Լ�ˈ�T�l���
v �"H@��W��� �O���	�\�CJ+*hR<��_J&�	/`�/��b��� �?GR��AG�wqq��8a4���a��K���+ML0+��L�|I0�q�7(���8���;�h�u��(�=8(? p��ge�)��|6s<���z�6E4�|0�@����T�[NCtGJO{=F:ymӒ/�yE���-����8Xə�L�j�Y��{�a�f��M��,rms6Q5�8z��������G�@��v�ΰ3�k�0[(�-�1�w����.�� ��y�F�8�7n��d;�m W%��	��:�x��J�3R�ʱix�p��ӆ�x���|gH���Q��7����f�e�n�S[=����8G62~�_�dӚ���x��aXF��48��̻-�+��t�[��/�3�ah�+7�k��s?�FMX�����h=��bD:��zPp�qR>2>Oa�@�W��;α� �~���]&"�w��u�,G���Qz̑�o����yfߋ!��Ox���ǿ~'�=`��IT�3��L�md��c`B�#3�����fS�;�ӭҼw�!�<|���|�<��%~���u,c���U��g7#I���@Zw�ݙѧ%����OԤ"S,n����.�7��i��ͼ�u�Ia���Q<��
��tKE�ʱbJ}�Y^c��:�;�v�u>�#��+�����j���&�ܵꜨ�2ez�{KDL���(K�2�%�8�v��T[s�[S	�H����w����h7�}.}|_�d��x��M��S�����#�s�#���O`�ub��¥�!�v2B1I��ׇ	��@ũ��;�%v�x�Ӈb���ش?�JZ2�H�8@���'N�˗V'dN��?߄dH;�Fx����`�j��l��f4 �=Vld����$9V�L������^Cn=RS�<_݌�R����Ș�1P�S"���L xa��^�u�`E1!0D�7c!��`\�MJ��v�[�JaG�T��7�D���AU���X�S̡p�$ߪYU~2a�g�-�r���2xe�Kb}b�� RHE���G�1)!tB��AΝ�W��T<��u^7�$�^貦�����1�'�}���V�J2�Ci7��BQ�����7�r��