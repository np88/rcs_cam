XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����^P̦�(ж�a� �ԓ`!�C��kI���20���5���m�$��*�9��j�����h����lph	p���\�i�}$f��0��̅X��ҹ�<�o����(�3��O�{ �D>uk</�<%.����f��X�a�� ��M^$�]��ў�ӱ�Az��W��)ɗ�e��1]~�Fطe��HX����+���<N=T+�������?�P����4�iW����������~�Z.)��ux����|�2V)��4��Ӈ�]���#��YZ����U�(����q��q�ml�J~S�EO�+�晅�Cq�˖�)/<>��x����w��&;"m���y��5�*��J�Tu��l�A0��o:RX��,���Mşnb���W�/m)����=�W��E�t�J��C����Jì� V Q��`���A#GoG����gf{�:�\��V���sV)�uaw��y�R��R�j�4K�!��-���I��3&�H�7���7��2��ߐ�
v�F����2���l��w;%ؼ���9���c����U�`�X8/�*��c�R*q�k����zd<��6�����9e��i���z��c����jc�O��
�W:ۋA��h�����U�ʀ�ww�oqJuDԲm��%���D��I}������`!�^�����O��eBz
��*Zd�՛Ѹ;�n�u��bW��]��X?)��+U����������!�-4�=��(���_%��٘k��:XlxVHYEB    fa00    2030Cļ���7�y�8�w*�?�{�����V"0's��D���Z��v���j�˖I@��V`,]K���l�}�����[�h���nz�VO��'H.!�=W'j�2�ȎU��|iq3.+��s9?9��2�{21��� {�D^Y�Xx�,S5���<A��M�y����z�jl�;F�Y��Ç��6ڶ����V�[W�u-"���@��WI�S���ږn�/�X��f��v�gd[��0�|D�����W0s��!��Ooy8�(���T��`�!���D�ݳp�3�+�0 iQ�Y�.�w\_Z:�8y���tfY���q�9te��R����n�\���/]}��ע�5ӞdX���%��t�H
?7CGf��ݬ��4U���`�~�1�S��#��b��j쏯�G�+�D�M��y��h%ʤV��q�g:�����͌�;w�?�s�|��OA�zP�@}�di�L�m9�uv��!9����Rԁ�s�\�J�z�4����%���rj{5�������kt�X�!fjD(9pW��4�eRy�je��\��n���1ʉ7UT�i�$�wPo7��ѥ�X��hB�1�6�	��%�M����@�?���G�
���7�`��A�gп�����3�K�������(8_O���@Y����nt��_��)X��	3R�ٿ�lj�_�n
�$Ȓ�V �����P6��~�0�G����A� �X�_�*�}m����Ϳ��-X}�T"d!��,���)�x�(i�8)�n*��!WN6!	�_΅�ı�*%�1酎:��˺6��������t���^���Q���*k����{�4��y�
Tq@f��֙��1>��>-BY�R�f�l ��{e|�@;�#bJ���A
0Q�?�ʌ{�i����u[M�UU�Z����HK(�b"� Wݰ� �����,�ʪ]Jذe����[
~���͘k����z����:�rƪ{U�����DDŋ���}�Gu�b"�b$��~�=�a]�.6���u���Di8��h���3��7�����������dQ���޾�Őc����V��B�o�1UG��X�W^U;��� 	c�%oI�u�](z]�AR4��S��x��,��=@��S�o���ל4�V/9`� u�v]��[Lj(��l�/W�Rt�xY���d@�~�C�a�^8�
�j�F�	L�j˝S%���T����r����@gq��ݗB��)�z��o���cC��{P�.%2S�B���O	�s�ǰ���\X�A�����j���}D��Š	�[�k�\;���:I�����d��۾e�d&5��4�"���	�Ac���G�i��5XҽHz5����������M� �e[P��c8�DȰ���)[��G��w8.�m���A� K�����s�lu�n�m`NpZ o��o7��j8���rjBԗ^u&$��W�\�Q׋M��QIb@b�1�u�	r5?ZI���7l���,�j��f�nh�-�m��n�wPʒ땄5��ުw�z�y�`&ʛ�J�l��l����\a\6T��{��<�蘐xo�h���FU�����G(�(,<L�\.5��m[��5��LU�ߧg�pР%��Ÿh��x��?���\��R��̒�ڍ�1��C�	`Զ���Nt��gáϩ�O5�V��s5T~֓ǡ�j��!|+{R����')vU�)�%��4��92�s������՗�(GG`�-1(dUA���,ʡ\��8��B��0���A,B7����4l[�3������
�/����%����T�vQ8QY�l��}��#���{��k۸k�Z��*����Y��Ql{0=��_�^�3e,(d�=1cK6D����#P\[�ز�u]ČP�����b��uƋ{��H� �ӯ�՟�nA�`G�����,9;��;HUG{��,���O��-{Y2z=7����cbA<+cBIS��U����ʓ\�;dJ�okNY��x��t:b�B7���Ts`����v�����![���/��|�vX�43���)w$f~�`\�ST9qۮ]�s��	��y��H���$���͓߱�w��#�JdK��
*2>^�d��S����Yެ�$�ǻ�1:�@)%Ã��>�!�:9)�!h����/��8�t��8��◭��C�'� ��n��y&n����\��~YT��?�dpӵ���k{l��y�xHЮ&z��Ρ:ec=�"+���M���|��g�].�D6;�g��h�o�c�{k�����x���bʪ��\ً��'�21�Y���GY�H�4M�X�E2���j���{�;l�� ��j��ܰ>|�.Bq2�7����g+���!Vu�x��T
d?����es�g�q&a��]��@ )�@���n�"�X�Ƌ:�ɖ��3�g깂C��
30�[k�5b�Y�F9҉TГ�K�Y(��*�}�ӱ��ߜ���Z~���~@�C�=�o
�
s��HC�hQ|�]%�A�e��q���V+S7�`�<��,e (f��ΐ��8d>
�i������(׶/;1:@,�/���T�K�t/z����f�ٕ��Jvns^<���Y# )5mզ�����T�Rѽ��!�N����`��Z���W����{[`��? &�,d_��J�4�H��~<��H�ْ��{0ݶ�F��Jw��ѵ�g^��<���HϤ;pH�Sm$�:)�(��D34�=(O�����S);5Ovt����~��
uIb��s��m�d��yX(�=k:�'�iYnC��>P�%����#��,�j�0n �,��������łD���N�=F8M�u��4����~zϜ
ځlt0}�x|ݓ&H��QL��̙l(\�t�HmZ�D�+7L�Z	��B�Q���`me��	�]�bo���0��q�@����w��w�4�BX���co� 9��&�����)��� ��!��q��B�6���7���CM8\���g��0iRN����ڐ�@�;p62K��z��ȼ"1�O��jӬ�&}�@�kf̵2�^MS���}jzY�g���쭨�I�.�X��ū�u%�'˩5�@�EǦ���/�z�S���u�����G�3Viv�u6C�и�R�Kf��ش����N����x�1�*`ꛂ�}��,Lm�2���--�4=�;b"n�g�H硝+iPGJ�����ؓ�
"���h�۝���9���
d�y]0��͵j��6�`�����EZ�`�BZl;E"(W����pKk<fD���q+�1�S�zwi��?�΢Ϡ���_����X�m�@��>�QpS�l�j��W���T���*�6q[>"�+���$Z�'�ѵ�m��4��{�a�^'��kE�7�P�p^!�~n%Ux��q���[d��A)*5��k�Wʳ1���Ԇ���� ?AU9.%B���#:e�l�w�T�u?=K/��P�ۯ>���;7Y�&�Q�te�-m.�lC��9v�}����@����-�m��j���Qp|�n�*��ˑ�}����A�[�}M�a��P�)�)\9R[�7Ǒ?{���VrT��CK!��-������]������&2Oj�h�f������9Fb�k��p���3 0��w��]H, �X6�հL\DyL�8��z�uĸ��&K��܁�5;�"�T��3˙`}	$��A ���d;L`Ao�$�U/'�41g��8Np �����ip8W�4�{��ɾ\�9+ZB��R1>D#{㲺�!b����k��� d٘����K�?�l-dm �����
Ȳ��X/sv[��vƚI
���Cw�%D��]>��N��a'�<�Ŏ6d!|�`�x���;�̣m��?�P�l� �E�hd�b�`m��>�\�_;�i=, Q����3�n�ſ�JR���e�4�u�c>~�x��?�ľ�ee�g7��!ˎl�OJ1���R�I'5�-��$���N~(�W=�Jz���~�x��F]��P|�f�f�	��]#��)Db<e@8�D�7޸�y�^� \����~k��#�TL�q;��(�%�А����ݦOy��q����HN�����_�ԜfS�@ã��O5�Fx���ݹ�W/v���#�IP$�e��Ien��h�>�H��Og)�H�s����q1}�J�~���i��|@����X�	s�1\:{0�VX��(���D����ـ��P��T�"t�e��RY�(�t�Ip��X�|q#c���p�o3�ؚuW��rG5D9� 7�{�>�6����_���ЅE|����յ?܄O2?�]0�!Skw]�e�'p`v*@������\�x�؃��^M�I0�ux4jus��9� m��.{��uͳ2�p�5��h?�&d�>>��p���&��1̸-/aBq���o"2��G�4����p�EZ ���N8t5�U�H�T�tOx2mEW9����F��+Y�6W}S�[��M�s@9a#�=���kv�8����x�5:?�9`�p4�,������f?a3	{���������q��Õ�c�G ��$�[;C��/����'äĈE�H����NPCoy�s�Ư��S.�,���k���j��yV?aFbႏ@;�����S��͌
Ǿ�5�3�2\���gUY�_�(l�M��b�S"ف��lP��$�+0hY��)��}h��Žte��ZF�c�U��ݞ��@�&��$�9�đ�>��y���RnV�2��jjHҷ�E���Cۃ�T���|�В��H��`j;�$a�wsɃ�nH���m���8�) p�����u�$yx�9_h	ۣj`��;�yqq&�,Buҳ׌aҾ@��2��.��#M��skYuHj�.�IR�R�r?y�#˩*�?eK��l� �0qm戌��F�K����ׅ����rbX�˟c�~Gu�+�� �'T,���J��cڎ�j��yF�L�ʩ:v��:,��;uX��_�-���)�T1A]�>�+T�3v�5��M��o7�(����FGɿp���qU��J�����cQ�^+�}$�-�㪊��Ki�XQ�n1K�]�������B`���7���;K�s�6e��NHX������kw�����j�1)	���<�U�f�q�GUW�/4�I��Yؐ��1��[�>��v��lW�X��"�k3r {�꯮���ݺ������Q�~C0��=|1�����K<�Lja���2cU����C'�De�^��9�%T��Yg>���_s�ʞv��ed�ή>
U�����fa��`�|����N~#>cfq呺w��)o�Qc�"�M�Pq�Hʏ�2u3f���&����Z�fy����x�(��Ϯ`����v���b(�)8��U �?G� M�e�_��ڢ���z��[ל���>��#��X��b EƇ�64��R<����UwLJ��ㆯ;5�0��}un�]��+9b#��\WR�'t��3� �h�b;>�ه�����Lz��gE�w�(�۪��g�x�j���+ؒ�  �-���<�4���s�z���v�k��sh_� 7��.��|=C�����> ��m���k�i���{��� �B#jqZ����y�Bu��| !�Z���P?Gu\+�#�g�!�1�|��~��G3Z�V��l�&1,�@u����2\7|`$�z7����%�e��Hu�zx&���P|V�C#�^��CJE;&��NʼZ�a	x)��5��vJ�&�q__�����K��e4�'
�޷��a�4.L|#���QGk|�a�c�t��s��@{�L`=�p�|��P�?��m蝢��4kT�i/����$J�Ufƌ#>{GDIu�)��+2�4�]-0M}�:��ݼ�|x��.�J�����"PE��y�(��v^VcZ#����i�����T;	�>����Q�-}b���"O�� /�_��4z�37wH��2\^#V��pP�ĵK�:������|?�Q���㺨?���hȸ��¢��=D�E�ĕ� n�߫�^���ig��%���g�����7��.��CÍ�Z�buZL@`<����0[7g�HId�鹟����r�����׊�k.���=�ܒk.t�Ĝwk�f'f��;u����Q�6*�X��G<R�	�X�@7��M`+�ɛ��n�����K�q�!Mٴ�<V���GA24��z+EXt��~�_�?�˒��o$��^��3���-R�{S��"Q2��D��h��;�w!�5$��O-M�_ъ�R���c�%r�p:�i�� ���(%����N��O���5�o4�_����s���*�t@!�+�U�J㼙J��c|��3�k��u;!ޛ��qk��6���8��tGf:m�F X
��:w֏-;Qkby�7�5:��)��꠮+o�w,;�
x��x�.kny��g��'�m�(Z{�}w������QR�>�wp�J�c��,�@���Y���L�h��m&�}S�7�Ѹ|�[�>߶�Y�Y�-��0��í}(|!d݌]C(�쥇��k�LQ~����
l�	Bg��_�$k����������N��=�ed'C\P��hzE��%�& ���C��~�*�N ��$H�I0xsC�!4R㜲������p'dG��i��i�����z�GԦ��ҙ�Ŭ�Kq�n�`�s*L����N�\n�r+1zl�^P� Y�u{O[����-���	�B���#�[I�Ά�Q[m�裱)R#������5W)�g��Is#��ۃ4�.S������i�b	o����/���n�&�W�O'�i��]�DJ����U�p��2�Y���7?�,g�ݩ�
�$Y\�IlD�5���d��^���A�M��}[�dYzl���޳"�|Ú�y���O�c��bH}e��
B����G=Ӿb6%-fU)���ڻf���Q�Ȁ���Aܗ�W���V�10���&�83ڷ��
B���{����b��\��ZY�D`Q�����oЗ����l9�9���:2��++0�~�,�̴U$��2�����؎��EI�Ґ���=`KqI_@8�^+��۝C3%#�,�~�(Ү�,�����|k���Ô� ޢ�cE�7����� ��m1	� E���օ3��ڈ�]� #�����k '/l;/�F��2p���?(��9�E��g�hs��i�Y�_7QEV����u{��!��{��V���ع�o�r�_��C���7��bh��rA�eg$��Т�w2�DK�K�/���U�~ )�͒X3UcS��=�&���ꦣ��O�"˓��q
hF괝�#7�J �w#�� |�k���Slv��c*�9'�6��`x�G�#-w�z�3g����`�qt��c� vc�~6,S�QS��>P�.��Zǩ���aT�b<�_w�> E]P�݃�[��eݔj�J*���[�'͋	�
A�yq�/�'	csӐr{娨�*b.a{�;5�@�^5�~!�Ë�!``',{8���A=�2�z*�ZhR���>$���PZ>諷ɲ8����l��ѠV�-fN��k�����f(:��$	���y=��������
��Dg�A�-f��߹/�;��R�S.snd���28��a���7˯t�Fgs�F�E�`��H`�mX�eN���?�q��nsS���k|޼�("C�JZ^Ap� c��x|5�Lg4����N��~KMx��ձ�:��Z�s�c)��cʐe��G|;�wҰ`�,p�$�Ay��a��N���uTM_�G��|E2";��3w�h�da�{��|="�rU��X��D��'���1��g� 0X?:�@��g�ڏ�w�#d�fu�r��+u�Gt>F=���Y��ה��H���5�YMA��E�i}�a~�5���t�f��;�	8,W���1ʮ	�7�wh�� ��0.C^�IS�5Bm7�"A���l���<G*�'/;��v�or-��K5L��_��o�zz7y��X���]�����nס`�q�����S��;H�����e%>>���;��*�`	�[��HX���H>����^67W�q]��r���P�	���x*"m�Ul�"�#���9��ݔ`֟��gee:+XlxVHYEB    9620     d70�{�s�@�����Y�m~���3U5��qܷc���V^���͆��ֽ�/��4�~d���~���T=yH:��"��u+�w��r諗&�	���X�+,F9 ���p��<���ey]숽��mp�&i�H��3*�C�p��=FJ%�V��B���"K����uW����)���a�頒��0�I7�3i�3]�.���|�ʶ�_S��*O�����j���y�d���=j�X�+�,A�U��NT�ɐÃ�*��r�Q)ߗ�
��meH��<A$�� �oE�*`y��#�V�i�W��U3��93ةv<��E.�ɋ���g�[��	�NI]��G��ym'� 8&C0����mY�l�CI��ΠS���� 2�^^}�MM�1�:`���D�,O4rd':�G�H���3�*A�#���5�.�M>2����n %i�հ�]���PCT��`����Tq�*�si��,U�� ]'���&����n�n#�w�朩U�h̗�	&*� �֛m�VR��e��=��A��|�k�n��tm�hl��H�!����Y�nZ}�
��^��S2�D��#$��a������,0Ҏ�\)�'��
�|jR�#%�܁�=D"E���&�K��q�C�5F�A�]�j���ʒ�W�-���st���}u��Jq����M��/�e\[�ՋW���2n���G?I���ɗ���:[g�
Km;���7�5s�@@)6����-JǅtȎ?V��&Z�,St�ه������D5���[��l�����������uB�	��H�eֿ~�6h���V��3hK�t�u�i3����4`�I]F�VN{h����e��E�w����]P�g�I����wV%�!�rd�!���A�m����|�8Q\�����?H6���x@/ }�5=\����5�<��*"���+f.L�@��۫�V���J�y `��%�s �&���8@`C��B� ��b��؍��y�j�QA��+����Oz`�ٹ�.�z)��q��(�B������=�z��2;҄%��L���U�y��C=53���@�	۴�j�;�[޳ gO�v��ե�d�)��f�yR �x9>FU�o���Ą[��qV����Þ;|2q��4���C�� �~SQ�F�+ɰ^O����=^}xSE�)��E&�=$�^�TC���p(0���U"\Wr�B0�u���4sGa���;q���<�]���"�~����I�$8�b��6L�XL3"+��V�lT��5?4���f/��sŽ��r�4\ӡ���w��:b��g�)�w�":��]�˝��>1E��G=��䪩���'&���[b�������m�N�$C3R�n���V���<�\�԰o�?��R?��B��H��C����EiY�ݻ�3������y�f<Xh
��hO�{��K|,H������>��Aa�m|�R�/p��\�,�//׬>�yĚ]����DbM/��(������r\M�������g1���m�����6�V���M~jT�k�՘���`
'8q�R�u�'��m1C�;s�zceeL�bɺ�t�~�~Kϝ%�oϝ�}J���x��"@��Zcqp׽�<R�z�=���]�r���nH�v��kdh�x�0]t�A1�
d��1.��ߒ���L�Io��\��l�,��ӽ��o�t�Ě��| n-ZJ�z7���?W��ܴ��[����4�0~�XS�D��@-ݫ�W�V|T�ܦ�"�T���2�p��M�5�'��v���UoK��K�]���|��ɗ��]Ш]��H�	{��~��x]�zƇҺ�3�]�I�i����"�����?�Q_B5V*L=�3j��2xL���,k���O଑�-HԆ�Z�;�{�E�ˡdrQ�8��S�9��?�8��{$��%&��))�:Ƙ���J["���i�]k��������ܤ�b���"���g׊�4<��a�g�z���k�@N7-H9����KP�be�\j֦;�:'��:7$kT�s�w�NN�P��l9���K^�����Ouブ�p�7xR�Yď�&���&D�^���'8UV�Q��v�)�)::��$�Ka�a���CP�h5p�x��y����?���sU����=�շ�@i�&��Ɗ?��׺�n��B��>��o�Y��r�{C�9��wK�z-~/TNW�ځ�+�8���_���q��N���q�)h�A�"-���l�~��oʟ�jOu��"�%Z{�^f&�_m�jю;�gM�����ZKֵ����/��  �=n(n��0͂W�"��&ܐ�&_ܜ_�?���~���y+f+y�=��׎�oKzyY`U�j5F��LpMU�UC�t�M
��oC�c0Ů��ߩ+~b�11�n~]���˅:��Y���׳���wnj��������zj���8�bK�~��$���m��>��Y�h^Y%JѰ�F�����1=�k)�VUى�H�6Uk�b&�!�b�̱y˖�D=�U��z�}Y�Kf�a�W<Tm*�3�!'�ɂ��։]���&�֢7	U3'����:;� 9f�4��Ć7%�j����I~-6c���û��pے��n1Z�3`8_��uh����[V��R�V%ˮ��>�4�w��nڡ\��"��:�a�����y���&	�,�j:H���a��E�k�S�7�B��I�|��c��R?*IxahG�WC�#Q�|21�{�m��m|A�֣W�R��s!�3�O1���|GfJ�`4ě�}�;a}�k���N;�(�]�Q�G��3��l���)�,�pg$}[�� {��q`���#g�������`�[P�p�='#R�fa�dkO23�sO�!+b>�����'�?�Mf�1`i�����(�₋Gmؙ���o{ԃ.�QkJm����/:OΒ?�ʥ[G{�<��%T�7�"�t���'�NM7��\_ڶF�k�S���G�&�Ⱥ�]�,:�N�\'M��	��,��{v��ܻR�;۱�<ƾ%U:�Α<>m�s��ww�����<�a �=�~��������p�\�\E��G[�l��r\#
��R*�8}L�5����96���$��!�A9h��1y��������)���	��h@�q�r�� 	*]��[��^�x�V�%��~���YW���l"��*�"�:'.3�nxxX�Er�v�B��&�����s]Vj����H�Ͳ$�?�d��?:�{9�+��R{mWo�kf���*gDe4u项92u�����κR*_j���NU>�ǅ�ίE�!/�_F���2�����J� n^���ĕ��p)=�I�fYA�V���ti\��n���*�]U#_��h>�?���@�f�.l+��*LU