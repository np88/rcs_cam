XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���������PX��)��x�7�U�V���XSo�H�294����ҳ�t �Zh*��W���g�N"�3}?ę9O <E�Kr�5 �z�Xg�R���(n\��G��,��U21����/S	p��&���=p�F��F�M`����:���Bī����e�lm�7ȍ�u�u�*Ē�`�����kt�
`C�Jz��c`��Y��7�8�k��� �l!���@W���Q��R{l��=7i���è|z�l���eg�\�iv��$�c�m�O �»`�f�ˊ��B?т�o�� u�j\+W��4Ӟ�Q�֊�K�+���+�8�r��	n:�W@6X��dIo�DC�{bx��q<�^���g[UE�F.�ռ}��W����E��z�H���o)A�0��Z�iD���Gx�b�'r�G9A*��d$UH�1�Z�x��z��<`B�vA��hqp�E�yJF�a�oc�B�d�)�����s��3�z�[�6��
������F-=	ji_�󜔿��qs����0'��裈��mab�����)�LlBZ&l	U,�71�Mn��y\�.�K~s�u�7�o��d����O�`�e[m�$�p�������fh8(����^jAW�`±"_��)Z;�� M�x�Y�g�����K@[��ge���j�[��J0�Q�FRp�<W��|�	�Z:3�p�(&���s��D%�� ��\�)A1�qI5ͅ^Z~H`����B ���Μj�T(F��N�CUi�xXlxVHYEB    6867    1150��5b����X��?,��x�מ],�eupE�u@|y�U����� f%�
aB�f0�8(�g�d��=��*_�R�J�u(`=w=�g�:�F�@�7�P�y?�<\�,�jŴ->x�[P��8���c�=FY�C&k@翥��<j�Ek�q#q���5*��P/��o��Rs�:��7&;�ЅU�28Z/#!ƐT������ڊw�˥��J^��#,�P�6�9�Q�"�}���̠�2��B��-.��O�1YT�������:��D�^��%�f��0m�uW��DtU�'&�g���A��R#�ނa��Y�'���`|H�G]���
��}�l ]�n�r��D`���*�q#��{Z��FA'�b��+�R�/˧~"���)a����^d���W�#�{���x�|�*f�l���NgR��fg�zGȲ��Y�*�$�vs���h��T?J=l]�.�!��յ�l�-4"T��u}��]oс�c�!BIV��sz%������f2?����{"O�ן,��֪��\�i��C+�Y.h���/@x��)��\��:9�
�d@��"�v	�Y6;�AL�(_J���i?\�6oQ�Y	��Ϭ}�3z�X�T��O1x�!�r�Ͳ�!���\
!�%�N���SLt4t�}�8�a��϶3��?�9K�T��6"ܧp���S<J�s@s}е�j�0CLd�i�UP���°Ǆ:�O,��/Ĩ��9�����_f�����.U�f?���~�#WT����i��<�H�� �ȷ��}�RP��.8����Z�kFD�6����ų~��*�8�yZ��Z*���SY�ok..[E�:5U��.���<J��75凢�`d�{RCR��\�9��H�~�@�e2r{��5��``�(yA���CT*���H�Nxbi}~?�rw�K_b�r���@	��VY��A$�U��h�f��J�	��u��YT$�/�mW���4	��(�*.V�kv�F������E/�Dݍ��Y\rW��,ȱ��iK�q;G����[G�y�����ҽ��9�]T�������(5\��C�W�x�\:�=�ZQ����ׯA���N��^v���B~�������������c�(2��wǇ~1<*��#\����Gm�Y�P:hWf��5�rr�� �G��G]�L�z	\�yuG������lX���:�*���h)/�ns
3�H�C�L�J��8��-�9=��`z>a@�âpd�,uv-��vy�p�TMaoh�E�=1�+���Ym;��Ǭ�聹s�&0u���"N	%���W�9�+V�ߡc�,>A����}I�Q��R8$nW��fFŽ�pB7\� }ͬ�{�wP��*��y��;i5�<�.�ZB}3�e���6�|���FhF���/=~�XA�׿���&��#�h$���b�r���������s��kmٌ�6��x�h�ZS�@��i���sf���N�AGK�� U�{�;�)�`�q8�}�܂��b�T�
���UZT�1�vfu��
��Q��4/VYb>���aFa��!o�w���U+�������j���dC^Y�(��}��d��]��V�&�� q�j$5$@y�bV`���'k8ǩ�Q#����;|7YpYx��|��T��%� κ,��z�h�����[nq�eͻ]"���UՆ��~�	�y�Zz�[�[]����H��K�|��A[��G������O@�C<g�p�u��������Y<��Cg��P��)h�Q*�p�#��[x�9	(z3Nt���d�ލ��`ۏw=l]R��v�@��(�fl�:�4��X2ʥ��r�}�F5|C�M�*	o̚��Z&���"��OM��e:�����8��v~:�x1(	�� ��D���cr�m&/����Hؙ�y"�.A��a6g���I��F�w�2~�-ۃ���������f�8�+��(V80���' S/PO��v�4m�`�����QC���_�)����J(5�@9-��6K<��<��zP�� /RX����x{��+�lu��4=�\��2=Eg���~�@ �G�U�2��s��6�JYFA;�J��w6	�%Uk��t�u1čĚ��ݨt������9h�P;G�)@D5W��v��wE2ح�	oO7�e ?2?�\9��݊`ˈ�׹h��0��q3���ĤGJֹ3�Um��VO�oI����Y�d�x��b��&"+/�3J�
/��EY<��ol����$|���G��	{%*���[l�:�
���U+s�-a=�߭l��ݭ�&?��\��i��g�4#�-3���\W4R���L�����V��|�����FX����R��*%�EwDx[�e��a~C�y7� ��f��g�	L`0r&�㸅B�f%�޸�Q�c��T2��[
���[�^}	��s9�4s�W ��8��"D�F�p��鯯����I	�^1h�{�x;�}���nH��L�1_����s�W�=I'P��G��lA�����[H��t�߈X�z�~p)C.��6��˥�RBn�"��/����ӳ
c��U$�I�PV>�?��#7"�$�pfH��H>���-ֽߢ��>m���D��K��N����G���O���z�9 ��gCaSG�G�ᶠ�	U�830����(�Sc-�-�v.Y,B��2���ˣ�ͽ+�:����k k'Yi��Jt�{ ���-���ܣJC�ÿ/��L�K�zEl�;U�3���t	��\�bK*�F]���Z�������p}�~�����6�"0�
f,�Rŷiܲ.�����4-f���-�ۼ^a߬0�j�x:MS�g釹��'X�(﮺0���( 7����^�e�U�D��K�t�_B�e�^%�~��{b�m�D���	;4�]X0:��I�����ebd�T�T�[ߋ����d���q�n�/�����YwG�Y�$�k���Ϸm�[�W�g�n��)Ƿd�*��}j�����M
*�_lT�!W�;���&!��}F���e1q�e&9!$�d�V>�ҭ[i�ex�c��-�`��.I�Do��E>�< ׈G��#:��Q�v�pG�Mb��VU�1WP�CW0�	ǫ�8�#�n���Q<X�qa=Ij�K˯(Xq�1r*��Eu��fc�|�F���i���v��ǐ��1�-^T�Ѵ�v������1���!����RE�!T
V�7��?�m(C�}���"��ǠO�E�Tt��;a�����NP�X������S�7�B��j(dg=�h��>���%���V	;8.��
tf\���k��Q�����Et�=�I�ό|c��mONC�ͷ�+�IF�2b�S�7�^8���-�\������}(x-h��9dAh�/`�)�����gƔ)�ο��+�*A��kH��!�^)9'�l0K���$"k�� ���4#��;��G'�.).��PMK`��Ro�I�O�#�~�����޻��8��/���BR6�(h�B����$~���0\ػ<�@nlv�u(�E�Rs7�<�틆�]0���t��)k� �D(�SA��fuZ��*�dE)����d	��Y�'K�j�s��|�ўcb{��:z>�8�4� 3�N�0��M��/�Y���[�ˤ	Ӯ��z���n^�`~�&.0zk��HN ]��1�
71�k�~����b��1d�_�x������Y.>����S���Yt֒tf�B�h2j_-��Y/�H����t�}���l�0դ�!LCs��"[�#�.�(R�m�ݭ��TX%�7��Erb`Bp�TA�a+��Џ���;�_1^�Xk����~
�^~ײ�y�y|�:���|`@�ճ���@�z��͵�y�M�N�B�o���+߃_/�C�U�e"D痪[�Ɛ@ ��p0_>���0�dI?U蘘� H2p�:������T�ǢW���5�G������o�D��S�߳$'%~�̐7��['J�Fd�}���;�Ռ�1$g�ǡU��n��k��8�A����ȑn#N���bDevꯃ������$��	�_�;�Ms[��*Yk�a���o8���Z�{d�9^�Hp����h�}�h�mL4��sGd2=��%nvw����!0S�L��N1Jxċm{>����{-� ��r��[�fw`��l>���%y�h��/�n=as�ף�xR�0��١�JXw� 8ke�*z��˽��ި����If��#�0���	S��?�l^�un�il3KIo�O��8co���(;gM��wC��x]��={�{�̶9?��`Y�N�-�7��6`À�m߯'�p���+n����C��4�Cdx�n� �I�z��|M"Җm�'����