XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��u�a��J%d�8hi�xű��,��&/)W�
�cT�1��d��a��ڊ�~=鍓��m�I��}��T�fe�lw���LA�I^�"�-�T��;��dh�V�O)����:���q�@`>O�34?άmi9�9X�_��h�/D�m�̎]�+S��V5���xG*�S��v�P2��1@�O��-�H��X���p@姕Ӣ+�Pt�.��i4�2�ϱ&�IV���`�*^���Œ����fKB���,���Gi�{}K�bX����/�8s��!L!t��)(�2�v�vƆ���<ܱ�O�Y��V32���~���&��wIB�/�ŀ �q�>�;��\yz�b=���g�u��#���R��c8;��1�\4�h��k��B�S�����~W3����,�&>�/Ci���Z.0ܿ4�|x"��u�"p̠\��W���Ȝ�����(�sJ_�Q����<�:Gm�jtO���I�'}�aT�&�y��#��2_b��
7��l�`021l��_����!�����Iݨ�ޕ��9���q�BFe4���_IbO_n6B���O3
�����/5�{�e7�mg+��7�y����5��G��
���<����;<�X8�J��X�#�^o.�8_Q��k���R��g�L �x��K?Z�)�"tB�sx�:9�BR�EJ�=7���V�.�{�=?|X��m�%P\��b��A���y���U.*�ԫ�<NZ!-�5l	zYH�4��� Sܴi�n��c�FC���d92XlxVHYEB    d6cf    1b30��r�d��uK��l,N�q��Vm�;l&>��~�������$	uƹy���`�?�nA�l�fG`���# �fKӻhܴ��U9��Ǵ4���9u�7\b��I|$C�>�;>�/G�Ỳ��{�����w�@�v���LG�^�#U�����Hv<^�0�G��6�<&E�ʺ���G�+G�J�����r�������Jr�vJi��9�o���y����|7���.[��=c;_��~�%��o̠t��<þ�MisF��xSx�(9�*g���%��,�ru�>}���Y�附4�Ԫ�`(�̫P��Dơ��I�5��[t �^��T�}N�.�ya
0���Ze�Ҿ�+���6W��͔!l��p{"�4�i�/���@Hz	@8̡�>�������#m�"��G2,]��A�nb�J֔��]���C���d��Q ��'�ڏ�qJǣ���"�WM��u܊�ޚ��?�6T�r(kQy �{���&��cY�]�=J�.���T�� �*m(]������`��Г+YY�=�Z��j����j��3�񞼔Qss2�u���p�[X�0������P���^�s?��܁�L0톳�ݮ����u��7���K��������^+�����#6W�^R&�Yb�^�E��ڑ�W���?tk��N�چ�E�Q�hk ��+x�%�d�(��0�� >�ħ�5��'7||�[?�F��6'�H�zZ+����,�8��e�V7��Dh�`��=?v7P���)��#�p��<����P�WYgs��1��`}����K�Bd�C�b?rN�N�����4-�~"_co���h�?o`���o@�Ȟ�\FE���	b9ɹBS��2	5Ǳj��ʌ���t{ofv���E��~x�.�of[+�3���ʎFM������%F&��9�v��v)ݺZf3�14c\Fټi\��3!P�B�n��16$^f34.�J��V��{��
�
S��^�k�N%�OM�d@wnSd��^;M�2���Sbu��isد#ǫ6H�8}��{��P���V�.B��ƱD)I�_\�����Qn�J���㓈t��K�I�H[�O�~{7�d��Tj)����� tmb8����b�%���1���#���-�ޓ�i��H��O�J�N����S10@sqYd.��#�ѕ�S-�t0�\9>r����~X"ر��{�;�F��|2�aR�o5��pFR�����$��t}r,3[�V�8�C0Ļ"`��3���a)	�<v�:(EnK��v�H��9Xd�����AO�Op�x,�\%�"�}�V���Æ�;�>�D��;���DWE�"Ljo��T32���r2��B��ȏD��s�����ϥvD�Đ�;�7�m��/��%l:�U����o2�Z��b���Xu�0�g�g�P�������ٕx`�')�;(�0X��43�;�=5�wHj:�m»M��Y�Z.0<�qc�|V���,P�Ѩh��
yL%S~�!0P��;N6�cV�(��E!?��ߧ�<ij��"�0��s�K��!����Z����	��W%z�R�&V�z<��_�@����n�1r[ym,�?
����+�{�d���0�7'(�U��j3�[C�¡�V�b^�HߋY�_���)k�bL��jeuղ[���]o�<�$�:�:�	P�;N�d�-��!����F�Խ]M*uNB�~b�sq!B�Ò�,�vVؿ��^ˢn%�TC��O�>
���Ձ���U�	�2�F9�t6��Cyyi6ӵ�k�c��7p�$z�m�Sk��t!k#��!-�e��Y�fK�/	�,����+h�D�||8.M�:2X�W�C;Dt��)H}��U̢�ril�Pj�N�vR{⇰\WuMקSh��t�YP�sMFD��RÛ ��l��p��~]O�t7��)k�Wz��J��ђ�7`�;�Y�p�YM����[
R������iS��nN�X����?����B~ʮ	�C��C_d[v�Pf0Kեe���%�kyԕ��D��v�p0�f�p�:_ee���>k��f�G����
w0�8�%hU�'������=�{���O@z0���?�c�:/��gC�����t�i���]��=��:f��
���;�k���y�V�z�V�-����3#�.�)!�0Y(�}5��0q �M����"ݽ��&��N��%_������/�:�a���$�ܒ�ӑ]nm��L�5X�؏{>iĩ���_t�5;��D��� :D�:�]�!�؃�)=�p���b7���:�q"v
��.�'�'�GZ}#WO�s��_v�1&�%C;Bvg�+]A�,�1���,᷎� і�}`��O�:���ԗ�Wq�H�_t��,푫��C4W��/�?;�"����vn��v�9G���n����>�p�jk���-�
o�(�Փ%³.!e8��;q⃙;�{S>�D�p��&@�Zr�~��K�?�$�,��B3� ڛxAN�����.��&����_*��$���k����`<���Ξ0gR����':�=}ի<&��E��d�v�C��&uh�l>A���I�O��߾Nv' @���c�b���Qsħ@q'�cR=�x,�"}�ߎh��7��р#�}Q��:�Y�q�Z�N�?�k����N������N�	��T0D�<���o��f�P}8f0;�-���ę܋U�� 44g-�}'��*�;<P�9��S&YV����!�����Hg�8�ɵR��2�0�&h�@�ž�Gsmo�����YA`�#�i�(���p&o���
���M����}=����հ�x�t݀Ox��%�׽\+A&A��"���X�Bd���0�F��}�0Z�N�#�Iu�[��V*v�2Qw��G��k;c|9H�"��\R�<��˂-�N�fzd�e�bzj�s�)���v�i%�5�q^��C������^d@_��ddrV����Yt���ݩM�!��P殇��F1�QY�� @GV�d�8�{�[�wҌ��3Q�����������m�S��ugf�ݪ�Ӟ&]�*���T����'I�8{5��L�-d=:�X`�����S����*��C�Ve���� �
�H��6��.�牄/;T�f��f���y�0�piʼ��{�J9����Z�;�"
��o�SCpϬ)�4�_��E�α�#7Z�ͯ���`�;O:��LSf.j���F\r��:vLOG�z�s/k�.���T��"-��$�*_�<}K�b���؝�vbak�n�뵘�L�lT���RR�M����q��3��+2M�K��(X��r^��9��u�ީ\*9�	���ŭ�k�k�Rg���9����H����n�"���=�o}'��ܪ���8���dc�\�v��/�ej������o��~t
1�y���,�n�m�R�)?�۴$�v3⯩=��>��OJS��Qu$~���]�� I7�����~�4��nX/��U�R�n�&��c�5٠���CeR�m��D�t@�ӒB����bɊ��ޗ�'lCҭ�-�E�b+rgc�92oI���E7dh	 p8B�5o�"��:�#��i?]au��	#Vw�W%(G�;�{ �oыX��U�jA���ٽ�]���w)>}�nM�5�>/qG���I�w��)�iT��nz��Ԏj��s��@��l�I�zq�"
��c��tX���~�6�!2��V�%��^����y��ʉ�G|�Pj�u�TA�����S 6I�L>�gc�i�\Ru�}���F��=۱�`R;�U�1��QED�o~�����%m�֧�m���hSХq^��L7�;��� ���ؽ\��(� �k��e����U���o��+�6���Bv,�ݮUNxC�pC��򎛘LF�g�
\���J�V�R0+}��D�a��S���	K�RU�M�n��S�7��K��,�`���~Q��;�;��W+���B�5���A�[��r��H�A*Y]����ż�ӸfR��-��!��<
��.R��I:pw���yh���/*4��#�W
��Q� �D.�Rp	��қ$.���E�I%�da�}�9��r�ȭY����.�~w����/���\��#���q�%��Ze/�'Y��laB%0�X\!SM���-z����A�f��mVC�9��	�����s:��. ���6B����yS�B�~ݍ�u���P[A��o����ź�
�*���<�";�z�}l�g��Fս+(�Aးm=y4ʃ���|l�A@2�}0�2�$�������9�	�1P��h�\���VD��#]6����YY�(,��i��P:�*J�L|�G��I�.ry'�Ϣ_64f��6�rB��֎�*K��E��N��Jf�"nLʫ���Ax���%���'$�WNB�sD��D,��i.�D������k�.�|�=��Za:�YB�+Yo�G�^읩?e)6�`,J)��xȆ6�Ir��5r��a*�i�����`�|J�'�Ҟ�]�
��K/Spz�4����k��`�\|��[�Jp��mĲX>
NR�;�#�����sjPjYɀ"A�ꏗp��NY[�������˸�߽�Z�J��>:��֋q���$_>�6�dy��.Gh��ˇJg��'C�օ)��+$=��T�a��:=��&�&�#�%�>]�x��d��?�Qre�I98 ��:88�}�/;�
�/w������6�%��x�)xgKB��ܿ�������8>֛�X�
D@���YP~8@���nkd
9x��$T�̀j���OЄY.=R�.�j\� �:.Ó�`��p��*�K��~�R2uq��}�n�����4�ꐱH~9��KGj�����b�#,$�R���\�^^ō8�qs5�QN����/�v`���pUс������N=�rS!�x�*Ɔ}���>�}��U��]�Q���z�gK�ShyP���b��w�e)�}:��u��Mu4afq�0uؗ*�o#d/�&�����9,�o��ڕ
�P��Mo�T��9�11�iU`�u+���ذ��N���Lf�=Ԟ�%5�v�SA�5FW[������bTm�W�҉S��\�Z���2�Pf��@Jf�N�v�';�M�l%�n�I�/����/��[s̈́Ӳ�����HXᬃ�.��K*�Q�D�z��WF�J�኉j{Y�E��?� ewnH��v�$\�o�e/`��o#�j����x��5ol�AyP�o��h
,Dݙt���B6�=�ɝn��[�+5�m'�@̄sK��ޘ����̍�O#�Xܩ���k���B�h�y<]��m�����SY����/��4?���/m�c�<��Mnp�TI����j�ع���(d:)�>̹���0�R�n<p�K\�&�j���m᷹\��V����/� �Y(Kg���)�xKb�N��fB�K��.�=������.�.���>lDx#_b@�WD�Q;9Ee�J���tk�Up�Dˠ����aѲ�	E��3���ph`���=�Z� �x>�[)��Ž�&�(�i,SL������U돥n����q�������YC*ؗm&{��2�x;0s#�|ߠ�Il�B�fGUF�Y�o�˨y�.�d�o��x�[�8�آ>�F7�b�`� uC :�cw\4C��Ibo�N�U�c`�U��!7�8�qe%�����Ni�g�y{��r�F�k�C2�5 ���_異�7k�t�ˑ~��%��JT{:�)����� ��=��5�N�M§�C/^ØJҝ�,NK3��� "I�vj
�r���<:yq"�l<Nۢ='�
��y��*���݇��g!E�F��E����-��`|U��8"SS}�P��9��}���^����ZH\#Ӈ���*���������Y�J�St�`��H@�D�,�?�Uuk�����c��)k&6e�))��qs"Ǌ�NQKY��Q��B��Uy�d/=�N��xtFq�� 97�,2s�Yݍ�B�nl��y�U�������Ȫ���S���DzIЂ�3��1��aKû�$>�P��oj�����@�����!KB�t��gZRe�T��F(�ꔾaű%���F�X_UB9��}�\� K��\�ćmR��X8�{�>;����\Q=����^CkI/d�@YO��EL�.D��VWZ4����:�>���9;���F�V>`(�����|�9�ل���@�&����%�[��p�r�Y�8�6�V�t?+x���X�ȱ��x�>���p�7��	3�}i8��;���1�{ۈ�hIv̫�����_m��|�����[��
���vn�)4S�v��Z�,{d�#�ڑ�ٲ��=	9,S��͝�F��/I�p��R�x=�N��1u_	g���T�<k�	�L�y���.߰s��b���B��-�:�p!�Ǎ�s#(��"��Y�vǨu�Mх���-�Gg��<���A���f#��Ol�:\t��N�<��Z.%��a�hM�_n�ʫ���8{C��ue]�ׅ��k=W�(�gϧ�:�9Iq��ϣ������5K��_��>?(���ұJ�0ma�m>�	 �I �����Hj�Ǐ���h��lU!z�~ɒ��Y��-݇8�H���|��S��k�l��"�7&�4�<�p��m�Ogά �@�ܞ��
�� }�x)�^�?���u��+��c�Y+HU���&?+
��/��X |ַ�݀D�+γ�u��#y$:�D��w�y��x0�`�0��)�����|[�dg���z_�Xq�U�i�e�B�d�j��]x���:;���F�i57:��Q.*��.#RS���d�T��
�����l�F�(��P>�Y/p{^*�F�@ ��u�F5%��w�D2;Җ�K�7Co�>"g~$CȄC�
0��Y�\�A�h�G�RѶy