XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��o�:�>�g0�a"�`���m��x��O/^>��Ͻ'�#�2��#��W�YR���Z����a��S�J}�-��a���CN՛K���h컦U�k�W%�������Ȫ�Hs�4��$��ťv��[��#��`�z�������
��ZgJ�H��ì:x��}xV'*�^l���PMx�|�dI��I������Yb���k�"Wޑ�B(����vŜo�㟤sg/5
S�#|&3V���R���l"�]Rk��1�'8P_H��B\�;�\���V�Ukp&S�틠Ո�U�������<�s�(�B�^�m�(����0ב�y�Б�;��!���֠%k���[z!zNE࿲��i�֗�I����i���������ٵ��n���8�:+I��Ud�����0NJ���6U'�w[Sn�d1�#{ ڋ�&��t�7�Kvj�G1d| 	Q�\��B�����a��~��,�Enq�d�i�.<|�T��^�k�z��i������<|�Wɨ�"ߺ�X��5!g�&Q�U�<?
�PS�BC�z�}�D�FM=޹��)�Ɪ��^�;��e�D�|unڅ�E��?_�NW�g���;�Q'�לS���P]�8y�;��uo��߻p릶y% ����F�l�)��C��\(E���]�
�����,	�I/�ʨ�`�JRN�+��&`�R��z�=1�rQî�ڼ�4��N\3������;�"<WK^"�[E^���P�xx�h����]`,
��V�}��6�XlxVHYEB    fa00    2470����!���e���Z p�n�w�-�5�3dm%�����4��42��=I��(��S!��^�{�\�Eq`�K�F�0��N�cM�ia�����5����,,��6��b��=���)�-�z���m�"Kr�ޚ�|�֪��v�K�L
��,�0�*�S~g�J"N�
=?�F��%��K���y�Kj3�12i�ݥD�N%�\��0�r>���E�Q=��ݿ��L��ym�l�`{D�O�;s��MpT7�Tf'#n�!��'�o\ȹg���8�6��)���P�gv�\�ӐIVB!�}滄�gpŇ��'ഛ4��ņ��=���`FSf� `�p>�lM�t'�#�$Z-����CM�<D���_S�c�qx�~�6��e}��x�$��r�	�j���R઎�5��C����7���7�F\�&zY0x��5�-��o�G��'���M=��\"�dF�T��뇉"��q�W��\�B��6�vEe��Z��r��t��0�=�0�X�>�B�#9y�=T�8���|�;X��3x�}�O�Yh��ڎ���ἉP����[�0{40�>*%��-7T#�3qu9c����=[>�v���g�{H4�G1���2Q��n"�#'OI���Z��mb�"�>\�خ6��L$\�T���4-�]�B��=%����=�����pL�%�!�zU�T%�e�D=�Y��ޑN*��I]{�ݙ�p|��0b��p�1M{���ؙV�^��bg�#�޸�f��l�v+0��r%�c���a,�i��b�V�<�;�F<ij�Y�K]͟74���|"��g{[����>�9!�8:r:� g��S��ӏ����q�,K�T��ahƳy=�>����I�sb�I���5�֣A��$	"lE��y�&�S{��<��#��C�U����٠������F4��@��.T��p=.55�L�/<��x|?T:9�L1�ː�j�H�n�b��x��@٥�X�h�m(��"ՌÀz�P���)�m�*�2�f� (xP��!�n9晉4,�����AUQ�@�Oً>]�Qy�ar�8H�hˎ���`
b���P�� ��]���0��Z9��[����^�w��3�8Q?�w�!|1{,�-�E��\�3��ȏd��ģ�_�a�ey�#mF��W�W�hѵ_'ɡ�f�����j�y�ڒ|��f�5�	�x�Y>�~�<�����<'��� ��M!�D"����,n���M�ʷZ/\�%��FO��2NG����T���Cdn��#��/*Z�c�,��{�Lc��� �vI���:I#0~�ﾅGIX�K�s�ee�(Q�'t���ɻǎM�l	�r�1� ��1�);Vs�7�8�`�HB����R�ˠ��L�u�"|I��[-d~�h�H<`#�J8�Ѥ�K],���3����k��|���?�S6�]R>�B�@�w��Iއ]'(�a?QY�G8n��yl*�1BǤ�Sײ����S��#p~�j�z�B<�7����(p�*��r��E�yD�+/X[�~�ij�]���WM|���yv���Fb��_�0#��wڤ�����Ӵ�W�hK):9R{�Bmg��O�t!��s��ʏ8�-"v�l2���E��H���r�g娕a�;��_��vf�W5ѩq�WdSR�sn�����3E��UH������>�-���/� T�9n�U����Y7�f�'F^���	���.O���|���|L���el��2�eS����Rx�w����T
�\�J)FA����p,�kqm& ��dU.��t�G�����;�ke�:�6���7�J<���7R���r+(�}�36~� ��m˰��<WH-�2���i�Z>VX�SK��0?aH���ʁ�7ޑؽl�(���]�݂�3��)�W��<�� �^�[����U��~�������W��	~��t��ۭ��Ë~�r"Bۥ����Uv��Y�!��a��a;W��J�}�)���u).c�m�x�e���8S*�*���x��b��L�����f-:%������O���ý[�	��`�Pu�}�Py�k
�����<9@��*�dO�2�=J8y�Z��2Mn�Ɩ���JU�橭 ȣ��q_@M`爉������7M17ɒ�f�)������6�d�tY�P��gN߅�)��?��H-���>�9��kL�!��ǂ; �j�qǀ��мŕ	9�rl���m�p`� S��Ş�8�UWm��T���Nc�pY� J����xYA�^@��ՋW��ё��PLt��	���� �äH��,[r����ۅF$��M���T_G���kLm:���ǔ�]�hI���4�9cI�D'�Afs���X�����k��&�g�8�c/n(�Чux��]!X֦J���m �'���<j���o�� _n��Ť������;g/[���؛���gB�C�{�K��,�]`�(�WOn���^C^d=_,
���,o��A�|Cѐ��7����#ٴvI��16k���>�$�uU��e@p*x)3u�X�^}8��oLE�0�s�(a���`¨���P�8��@����U��E�=�OҒ��O�@���V㞶%�U�D�� l�s�)�8�s����#�tDb}��#���汥-�)�`� �#�o�@�`�Mf��o��'L2��n���P5�M�ܷG� ?�vø?m�i�ڔ(���<u�����Z�-S��h��$@�'6�p��(:x�P�:cU(�,Y�A�s��B���e�Q᜙	�*_���+Z��#ߧ�)t�}��<��灨����a�F9���1���sv1�|II�C�φ?�[��k���~��D�EN����"{d�x)8T��g ;8��6~��I��������	a���>٭R��3w5�һzs9)T{��@.Xa�!)9�o��_���4PJ�*u�a��`�drY=[?����/�3�փ.����G�痏1F���ZQ����5d����&v����3��Ii�*Ğb��I<~�C�m�K𶧀=VGD	���[����yʅ�7��Z��ڸH�>�����}ng���{���ռ�p8���C�X�:y|����rH�2/�ן�3�H�"`S�j�����w3��*9)E�(�Xz�uo�V^(
����[P\3�"\���3�F��d�)[�������V�̎Ћ�(�6�nJ���� z���X�
?"�66;��7�`��n��;�
�T��b�������
�}e�C���L�&a'��'���lEG��r�I�X�P�x�gq�F\�c�ďK N��\)[�1�� �Ӈ�6�b�`��'����WDz��GC�X�._Ù�����Ild'�@����&,��j�a�?	�	aF�h!�7�G+���2�Wh�|s��0/�D?��ĸ���V<J������A?א���Y��P�4}����C�*A�,�{�܍P�g�����6.�;��ُ��q���ʼJ���;I����5�(I��~��>Ǔ������(=U�2���W�Ad�z���c���q��9	�I�'�����3�(⑓���ȹ��f��Xߎ�w����XAЖ�&����7�<beU_���o\։�ֵK�(}�A�1Y,�#�/ �?��)�Όy�e)/g����
��]h?'\#�n�B&��F��Wx��H^E*����n�pa���R�V�X~&6ߗ��S ���f��4̿��F���QP�p��N�]X�v�t���9R`�� w�n	r���U?��jEn�NPZ���v�_�z/��C|�.Θ	��k��+�v$�J�b��OR5Қ	�$�_��4� �	~�אie]t����vbI�^o�}z�.Z,���'�T�(�%�1�գ�?;��[���x/+?�����'y��/���~m[����% �j�r�Z �I��a��zHY����΅`�Í�����Ŭ�5������iY��*P�k	�R�'I��Q�#<��2�[��|�2^ ��\L����\\)2�r�@�Rj'b��*��k��/7�u,^�y/ ��T�h�M<T�(9�u �>N4#ZV4vz"$G҃�i����"�v�w���6�\k8Ani=B�g=���#�V�����NIxl�;U�4�0�c_Ҭ�z?T�5���v7�ߝL^�����3
;�������8]7�Ț�t.��}=���}B� ���RO�	Lm�%��f���+���<0Kxkn�^������R}i���FU��]�	y����&��Ls~1�fh*݃�BE\AoE
�C�ױ�f��Co��v�p}墇6����8�a�q��/=����Z[�JX�|n��T<���]j����R��di|@�f�Z��2�z�Kjwj��;{	�.�r�9�5����!e؉ʿʈOT����0T��#7��pˤ�<i���|�[�m��-��Y�iTzcۓ���(�9����\˹ڐn��E*nv�#��ρ_�yR�.	Ԫ�+��u��Ԯ��ӂ���p�0���+�s�k_]&:�+����l���rv�ج��&�xmm��6]b"�a�����s�q�`�I�7R5X0LJ����t��[z/x�g�đ�x����`�5��L�r�D���C�i&��1��ڐ���I��Y��h��oc�c�?26m1�S���-��M��b�E�
t��^�r��L�1���4���tj�����Tx�o�q�=�����mE���o6���k)U[ǤH�n�-�e�:����l ��7��,�z�����Y\TQm��S9�4�4U	����z��
J�6'�h��OA?5u$)97���e���{�}	�V3.am|�k���`T��X*�)u9L,�-��{�h{�PxK%0٭'pPV̭� 9{;}<�&V0���]�F�U�{[#�eT��5��!��°p�u8�:�@]3�-�ٜh㟨�!�܁!8��oUIi0N����9m��#���&M`�Vl�N���se'���US�7��.h�M�I��� �s�UM�(U�P=^p�bF���M3��K)[�wԄ��)o��>i�.�L�X��м0��J�ěd�Ql./J����Z�����]�����@
��k��p�ȫ8�`X��$d2�-�$�a3�Ԓ3� ��ҔQT���7�T���x�"�?;v�l�?c"�	���l�;�sv�&��-"r�Z-��#M��e�m)|�!�C 
�r��D&�����VK��N%�fkU੪f�c�kQ��R��w�*�-��병�s:�Z7�i�nɳ��D�1�r	��D0Q ؒ����7��Hb��e����בف�;4�	�,Gd΋T���^5�J�P�,y!3P��t/��_X�O��kB��b�(����QX/��J��j���򺚑�=�-���U�mw�@YI=�>�|F�6Y�.5�N`������+�z�PHD�;ɧ�]^a���o��pN�\�G���R�+5��&3
%=^����Մ�0�H�����e�a��K*� �JQ�Dfe�S��.LA��1E�GtPJ-���v͗8o��|��8�0����K{*zs�ۜ����d"q8�|{�He@;���B�7@��&��ϊ~`3�drf������p��ӈ��in�9 
m!��U,��	ޟp�m@�ˡ�x$��ĥ�d�3@�#S~5=������v����������Ҽ�b��]����	'w_�E�<��Цd��Ʈ ��?�X$���?�9B���z�n���=U��a,9�o�̓�|��t ���AG����&v�>�>u0��39Y!�LK�1��� e�0��:�cL�ŻO�90�xF�Q�olOg������,8�\�s�v�諄)q��mx�e�u,lz\��kjFBt�	N�A���N$���#Q���`0&��ؐ�<�kިs!��t���t��z����am ��y��j.���4�J��ܤ��pE�S����poً��2� �r�����!q�.U��g�36ǑЀv_���Q�f��'��&�l��IO�7쥾��;3�c�<b)�u�K���Ǚ:b�4�7#IGѥ�*��("�R���.p�$9*x�݅�w�D���,<(��x��5�u��W�s0]����H�2kn�N@bQ�#/�g�hcV}������b�8V݋�qN�/@�^z�:��i�f賩�;lN���rh���w�&���3�g<F��8�kk��~*���N6�P�,>�9��Uv�"�����*�1@ =�RD����l,&�s���a	�bq�q��Y�Zwg��jث�)�Z��],��|#����P�1��8���<�#�X������<F�hωk��C�/�S9��z��-oH��#��*Rq�j5Vr��<�Vsii^������ uɡ�n�%YgF�EG��l�����Ü��>���z����Y�� J%�R�6��2oM;c��
^S���A��Z�S"Yjxm�Z��z���
��S�`��*�e{L8��ɳ�ᖠ߶���{��>��2��ݠ ��u��>aE6���dR2$�ֹ��*���@nO:bЂ�}4�cg)�.�X�WN��ISԌI�Z)�_���O�9��\w�c�F�������D&�oT���~�,Z��7AX����@|������*�8-�����do�t����ݗE0\��(+Y��Q���g� $`��5c	�U�б�ͪ���>v����'�aX�`N� �	B�{���x #�9R������V��`v�V�zZ�]^Q��߭N��9�o疮�y�s�4��Jd~�\����;���-�>n�� _�9�Q��ʪ]O�4{�?�&X�Y-+��)�t�<S)��9&T�ʊ��d�k���h��61�ʏS��W��U|�m�ޞL_v�%���9��T�+�o�^�J��dV�����߷�)��K���4��F�:���<�7�HCdMU��� (P��-2�D��%�J��c�tIHHѫ$���; ��/tС�(\���~=jj@�M�%:^�2C=�����Ek�Va�rCq�$����y��eA�k��,D�Ѵ=��W�R���	b�)��\*��&0��spڴ4�m8�J|d%c�I��!.�׮&.h�����[u2 ��*�j.�����*��F��<_$���� �n��Ӻ�m	�������` ���/k��H��&�
*��,Μ��G�}�:DJ���4��t���J�O[i]������A6�$��3f�K%n��X4�Zͥκx��"�lF��-5��z��)�.���_�rG�k�{�@���ErN�cuwTx.&�K�@�}�Y6���$�G�]?L�	�6gseg H 쨒��1���i@�!��s�5����n�YH-[��᱅�%n�P\E��bPOm(\�_�i}����r�_X�*i=�Dq��/~Q�ȁ߰��K����l�6�L���]w�2�~�"J�ݖ�{�A��;>��!�4|�$%@��1�見�W��;%	��+�s��䥍�[O��k�|��\����x4}ҴM��.!��f6�l�m\/�O�2P���P���qN]�2Sx�<�r҅>��Q@��~f<?��B��̛�NaS����,����@�����)�l�Hc�w��͗Z��A=|��������?,+{��\�^C5$�uʴ����`oՃ�!`6���&����w�QjD�٤��?�gE���m'��Տm��u��Pi'0��V @}�p�m�Z�}���3��C�G����v�G��Ʌ �f���ٯ=[EE�By���gD��N}U
�A��Y��O�� c��D��2Jз ��U��;�V� ��ܶW:�V��/�f�J ��KE���C�l���8T^.ԗ�0lO��5�2�K�[�.��q����kf��u#��KC�
>4�@.)d6@R��R*;^��ʽ��6^9���^�)*����R����q�nM�ޚ��v۱�̹�x�K���4���/	�t�5����&����l{�ӻ;��%��� rU��=ԁ�ъG4R��%;�RL��@����2��By/ZY���6�W��8.f�u�0]6D�c�	�K�u:��E��4�ƃ��>aݮ��s}N���_����>S��G��棘�@��S�{������c�vK�'�G��\Ur�oFm���=_��s���D�L"��j$���К�x���F��g����3����l^�ne&��b[����.��PEB�=��+���1M��>�$;IdԜB5]i!�y.��������ǃf ���q�W��D����a�t0����';���;���|.J���vf(z�^fg͕_�]�"a�A,4n#3�6s���@�J���]6��yZGNj�.C� ��i#��r�URT8�osM*���h�-���sm� v}���#�^QO~�e��)�=�/��z,Mіܣ���cV�!��Ҙ�%�1br��=ݴ����F���S�,�1d�+��R@����e0�G7A��Y���]����na3�<3��+���Km�p�L\2�U�tB9��ؗ簘��Ѫ���u.k�Y�����`P����$�g�G����N���@I�JǤݔ�dz$�&h�mw~p˳J#_CIS�G���(����\,�t؃�ߣ6������h��i�LjK
$����ۍyb�}��[*�	
c/Q�%������_]�R-�_�jg���E�8*tǬT��/����S�&s���u��f�:,�#��qi񅥘M���{�c!yg&�I'$���94�����	^��v�=��J��r�I�� ������e�{=I�Q��|����`~�������A*$�?�-jE8#L�7�N���v��zV�����V#����6��<�Iklr��v\q>ˊ/��z�h$���$��ʀ6�mu�Y�_\��^����G�T ��H2]n˄�B:D�:�)�5��u޼VS�7|hȵ
 �qP�4��1_����`�C�$1���3���M�t�'�z��L����r�g�w��٢�#V`��������\͚��(���3|I��X���S�EH���l<����G���?��Hƞ`�Rp�<�[�[�/;W:��#����|A7�	�I�0XlxVHYEB    fa00    1b30�^���n�����ZG�W��qX�{Ћ�XꜦ���P��sL�6F�?���p/�u�kɷ�Z�.����G(�JĂ�*P6��S�Gݒ��Im�b��[JB����SZ6���&?�������uaZu��;*`�±���ë���e;�	���V/�*��:�t��縏ׁ����;ӜV��+�rB����@��H��7�{!�##�ld�-[ӐE@I�G�N�Z"��gK>�_g�x�	]$�},�i�sؠ��(}����9�󂨿�G8I���[�H~zoQ��i5�?��0*{C�7�	k�g��5g�*ƀ��%r0�����ت<c�V?���=�����Y+NS�4܎�h"8`� �7`�`���
���EQL^1ƺc�𗟀EJ��}$��Y��������|���2�8�4��bcYL�r�5?1���~KD�[	�r�N/L�(&}� cS@۴5m��j�S��> ���?���z�ŸL��!��]GUʗ9)��e%�U�`Ȓ��MS����,'#��Dñb7��ZJ�H_}�xO������7�S�v��A��Kb��b��SS�)�3�ԱQz��2Ky)�0�5�n��eӟy S��`�ͯd <��xZM[���$�Fk$?k#+�Bf@WE���-��S�����y%� ��d�e3ĚO
�U�}�z1לl�֞[��@b?1�������&0p���d�l�4!T�MH>��}��Ą��U����^��\��$)&0��,M�'�{~S�ng3��S�����`�e=1P�'/�_��P���tk6�:���I�[`/�k�ˑ5+>���O���sVJ���`��5��ń�сn�0��U����,�٬�=�:���u\�jxy�X0Um�$�g���W+�t�J���9����ݶVjY��j�$׎K	�ݪ�]h��5� U�8
8��+v�:0��ڇ��V�Bc�=}��8���J=��KU�76u�
�Y�=��4<�OJ�%VO{�~����f��/tc̀g��u�o;|1�_��
Ȁ���.��-afú!)SpNy����-�q��J0��>`ȮUp�����:4 (*��n5�&6�⌬4�TZ���*?8v�V$�tZ��+,�/�p�7�o\7�
����$t_�c��/p�x��?8�m���2K0ծ� D�pu;��%^SB(�ͫ+p�b��8��OE�l�=��J��&�L>+&"��ǣ��f���x���c1e��Hs��Bz_�*vI�|�:mRy��R�i�/��Krc��>�L�)��rF%�7��'���8m���f��-"Ԯ�uHu�UJ<�?������橺���J�V��2Լߤ�<B��X��8�FG�,+���|�������SrU��~��]�gm<SqGsA4	q#D19�;��ڤ(f�K=�w��e}����y��!0&�au��ө&xO� ��
ų��2�ѭ�,JR�̓�(���m�4-�/Qَp�I�l�j��߳y2\��ybOo��o<St�v��7N��ġ��Z�V7u����H�,U���7�& 8�e8��[�
Ը�y���9����)� ��&Jl4W��aW��&�@��T*U5E3��>�e%�\�'b�?�p����@����5L=d�N�h�k�� ҳ0 �TD�<�G}�_�"��&��� >�O8��;pL<z��{�pE�3e�Y������
��ծ�j�����u��/�F#�����dx0�����>B�n)�E�YW�)r��Jw�,�c4R\?&͝{,g 85+5[�h+ͅ�W�~���BZIst�l�LbPCgv�>��q�%PowC��d��*�;UR���m����_���ةp�͵���B�uG�/,����b9E/5�)y��Vq�?q
�Kq;�>��ڿ6��@S>툕�1���HSd9��'�@�����JU7�蹱pC��X
��xcc�������en�������|A�/'y�&���"%]k��аSS�϶H��8��j�s,�f�IZ�~�jpX�]v7<��j�����񴰟P������5����1�ȍ���ގ]B�"uyN�-O�.Y�"`�W��Cg�H�J�%����Y$W�(���7��rQ�a�Y/��A�q�F�F��-a�5���A�&n���q3�m���ր(a}9>M^+L
ۨ��~�ɫ��d���y7��b���xa6�wbB��?�fPg� ��p��OJ���<�L9������Z��Y��Z�I΋�B���e�wي��?W[� �`��^w��� :�n�4yD0�`�E��E�+���d��!�=�w]��}�Ղ�x�#����g&Pt�x�����Q��_1�P�7����4�;���Y�����Tw�O��VNj�e�@�zZђ�3x�y�Ug�T,��;h�9���xN���o�Jp�g�r���	8895�3�%�p�8~�`�v�tϰ$ߧ���˗��D�p�gΗy�J/�_$;���,%��7�s&�$��x�o�'o%�W�}���A�KC!ڷ��@D\Ќk1g��Ől��]��[O2K4����.5�ẏ��`��;�`J�>���6�T��z5�U�"g����6�$�u\�
r�7���$�8�Q[*�s������M(\����+�H���/�n�/B��&5��Es�]����ló������n���Q0k��4���9��;���n�F��/d:p����A�mֲ�ǁv��$Պ$;PV�\�9�G�����'D��(�sm�`4�,�!`�ހ�>��8�>�O��OdUa>7,�ӆØ{�z1��3�pp��X�nܧт���wg���*3%Y���u߀��0�7��,����%�c��*���K��Rw��J����1V+j��m�#�b���K+�S�����ː����ӹII`�ل�K|�?�OI!'��Șbzqӷ��w{���0�O`uLb%$��Dh�d�<W�N�׎��'�<V��O�=�zS˞Rk��)��j��#�	�����d��o������`��k>���ğd.��D��(2�_ĵ�ă�P'�=$}\�5 [������$�8���3$Gr���F�a	9��8
��
h�����_�WV�ϨК^��]����Z�1���'�%�X���j�� �o8_#�y#f%σ�1H��2`�����b>t�Wʻ�����cE�G�������%�|�3r�`�&����њ$L�6[U���ƸV?;#ĥT��E	q�r�U� �t��o���%?p��%[��Lǜ�#�;���Ӕ� le16E�ҭ]4C��?Tdj��|���������;�pNwdޝ�NW�!0�%����Ea�t��hܐK'��w�q��=P�����S��	��j�hŧ�J�c,S�K��Q$�!����
�Da��)��0����`6��V��x��J�1ƀ<C��ֈ�|T�!��ӛЄ���%^J-�^Vh��_��i��DV�-wV 3Ln���K�}|+M��p"� �L�]���+oWI5��=��9V5�(� -���(m�YV��\j�꼡�B���w���� �vX�=���f�#��r���W�n�_��y<Q�E߮�ë����V�(�96]Z��;0�M���L������� �Lg����u|�ٲ.r��Y׏Z��ӻB���ce�����%��jH��$�&K��΀R����`�2�QU��؜�i�s-���M#"��r�������R��]�@�b9�Ίg�mO���!��g8�9�Fk[�z��YZ]�a����`�R����)�_��H6�F��h9�J7���R�i��A�R`UuUN���o����O�a8�(�z]��L
��l�}"V�x���-�&�5���Z.��.�9� ���gAفoH�$����߷84���	�P�	�~*�1�u�Q3+kc��Ǭ�f(�}:Q������ۯ_��R���,.X��i<� Hk��ӕ���o��ː��B�\ٔ��Ƴ4;ZL���P�>`EVb����F��O�Ѿ���nͫ4YZ�=�ɨ��.�=�i�zˌЃL<�!kH�ͽx{wK�:Z�Jwn���
K�����r�A���HRO�.���)��a6�?�2뒏�ZN��#����m�O.`��sk�C�$�Co�0�w��{����IQ�ϳ�  �+X��N�a����.ʷ�_29���5%VK/�aF���5q�<C���4�mryMDԻ	���ޞp�/{�����B��:n'��Y�6�*僻F?D���/���E�,l��ψ�����i�毐��Y�_�7���&I8j%�+�4�].�ߺA�Z���tU��5G�ބ�B��6��MI�dk���-V�`��AU�t�X���B3U������*Z�:�C�~���gx���������Z��Rl�]$��i^��~ԯw��u�rX��C������p�A&a�\˗����>(��:${�
��ԩ{���-�Rľt�x�}=s7��n����U�EB�Ɲ�!�ɹ6��Wv�~��x� 
�Sn��6 �}-�����`�{p�2�b�/�BS���jzaT���׫\��JH��4���@�QǕ�Wۃ��o�������"Y��h�<jE(MBy�j"�A�����W�����M�Y��(��Xq[s��ph��w���y'�V��*u��w��6Z�G��W;"��U�e�ν�`�!T(�u����Z%1.�U�1���E[^��F�V�4�,����f+����T�Qq�	\��ߒQG�{����|��Y&�	ҥC���H�`E�Yƃ^�{Q��Sb[&/R��
�AQ��l������>F��|L�^����U���u3�k�M�Q?��H��8-���<�t��> �pu�����-5rN�X������Gx����^	N�@M�Qg���4=ѦK	� ��?D<EtJ�������v͈t���1���ؘ�ĵ�7�e�����T�tR�a%��(������+,ī�5���0T}���(H��Q�� �?nv�y����E/��@��CL_�ߑ��;�WLCz��y��C�V�Fn\ʟ��x;���v�T/Ŷ^�
l��>��\f��U��*=�?>M]��"�0���,��"8��ȭ^ 
E1M�{��*%��,�Z�N�!H�J>]�l�W�WHl��y�V1u=�`�u�T�2d�+7x?��>�uwF���IiD�/�o�:�)?�ٙ�e���kW�;�����%2KN�dF�߶�?;�e�E�����y�N׾��-n�d9����o�[�� ��=�.+L3������,�n���7r��==S����2���!fwK��xE��%���(B�\�:-մ�>��:lj=5o�f� ��gGI�!�U��5_e��#�@�8-U/�/��2�
���Ԁ�ݭ,sq�S>��w#��������R2ɣY��(��ݳ#����k:�C�ܙ�{��-���!6ü|�	i{x���,s��bc%�К)���S�W�6��o���N۴P<#u�����L0#�j��ʡ����8���WbK� }��(�r�GN[�ch;��r�K� (�aQ[�:�5s|u�=[�m
�Pa��M����d�k�TL��l� s���^�l�7�A��Bޗ6���X^5U�Q���:-<�A	�KI�)s��Wub+��S�SI���H	������~��ON���N���"��W{����A��Nַi���B<����4�Jr,i��\!����
� `|����?��>o#�ĉ�¸����<��Y�M6�<$��ѽ��|��ʎ�2M�lb72�b��� v������vEk�ru����W��c���Y;Y�R�_�0 9!�����R����Ў!��+w pNR��/C�?�6?��n�*}k���[:ԉF ��r��PS9ms�8��*�kT)�5�ޜ��e��qI���7��tn7gt���-gO�(�lȌu�!ʳ}DAvӢ��X�kĐ�2�ȾH����������`�E*x`t¾���[�D7e�\M�'1r?x�;��f�.�R��[�.���5:��g���S6QPcM�#�ϊ:���u�蜳�����,����Ң�٣��+��J��r�ũh<�N�W�z������-�ٜ��hKc �6W&lR�����Rz�i��Oq��-�}��w冼|3���x[�>�2��C�D���8�1F����E��wrcw��>�,��l�R���u��G����E$�U>h]Rt����r�Pa��� �âX�4��<?Q��'j=�T	W�䜶����n���ԚFN<�`R_��-f�&�mSg)���Wp�5?9.�	0�ԥ���;���C�"uU��p����Bhtc��^0�}?�����-�]��������Ra��k[�Tj�s�����?�\�<�ع��]�q�*m[��7�p�Ц�߲R�-tm��ǫ��!Ej��a��쉌���;_�em_��	�kTͬ��6^�ƕ�7��n �q9﹠h������@K�6{^�Bc�yҥ,� 
�X.����_���֐�r:��
ג��۹�|�߿����3 �F�B3���#W��6)��q�]��р�e.��Q>���p���<�K4r���Iԝ�Dg�Zo*j�Ͳ��OH9c;��9A��K�(� -w���Ev�i�Lʦ�d���V�,�1�G5���&��r#?\;�>�)hG�A�4���Z��ě9��������4��4�a�����M���av��O��ZS���˂����غ���� |�;pK���G�tJ��E��Km�|�Ƒ�j|Ӄ�T���-�8m�eYE�˺"l2���?���.��*qQ��N�XlxVHYEB    fa00    1950����(s��������B^�ΥGęHu�ً+�C�<��ܚ�z*�H�iZ6�=�y�-^�Q���4$����C �=��;�8C�p�9IKJ��*x
��6�E f���cn�XC����s��I�e�1�{U�&m�D�wD*6��$)�b�݇1y���KA�8�?��t{��TL|���i�Q{���h��]��p;4��-'�������n9��#Q�[ !��5q�kQs�o�sh2XCpB��ˉ�3�=\��ٶ��R��/ ��㧐lC�/�X�h���X�����B3b�6%o���ٜ���-�6��M��7�0,� �$��5 ��ĵk����;�#}����S��5���0�.S�t'�ɴ����,j��Y'�Nc�*�d�}�4�DQ,�'p >�>}]���啷~1 M��w�(�Ł���5��	ؙX9�L��"+��#�TO�W-�))�[�r+���!�< ?���J�����~4�GTT ��\���vc��Ә[|M�#ώI��f����#Q����}uj㋆_�^�*�Ks ��ʓUgv�}����p����� �v�.����&��Y{���v������?%c8>*6c�L;r���"veA�m�08u.����Va֑�?0�?i5��>�x����l��-G#Ok���x���zT}?0�q\bw�o4{�B5nsBD`���7(��R*3/K�=�V ��n?���K�#��I����|�b9`8����%K��9-L�ޡ�&�A�{WζoD˱�	�J�� �_�h@k`'�{�	$�K��Du'zcn2/|A��5�@V!�$���T�c�i�����s3xǄǵ�`�_.{�d���6r�:�ذ(i$�u�=��.�yt�����+ΧX�H�jYX�K2�c�4� m�a�;=b���u���+n"_ng���:�m7]\
�����B8yEc� y)�K��K�V�H�%d����^�t�z�ϥ�G�Ɵ~a�Z�P��,��=�O���J�$��6+"�t��h��V�3Wu����vd'��oʈ</߃3����5r*#yJ8�S�Wq����ÿX���?tS���(�	o��މ16`;�>�:�^���]���m��D$�P�2�CFQpA] {���!����B/g�1L�5�ףX��|=~�����nuy.�V�g7�*,�Ž5�GE����/5I�԰K�>�Ԋ�%z�l{	v�������;�|�!<^Mp��-�L�@�*����"�"%���J�=�rQ}�U2I�c'�k1�apr~��J(\��aY�A`1�`I^������OE.h [mWW�
;�La�A��Z%#Qx�{���r^+�w�e�ufQ��,��2�{KZ�c%��Lߥ�h ֆ�@:��ֻt��Ե�h�L
R�\���� �t�$B��^���+����ֈ>n�䉱�{��������C�6b����%��1��w���b��3�?��%M�D�4�a;	��������X�秪�%��^��������;�4[D��\���8���/O��!K����t��"`�@����RQ���L��r �P#��$6�m1໦�U6ꙭ"<�A��{}�޾V铞�	S4[��牲�����l���֡#�� ���*�R)U�D~���s�Yoy�b���4�;Ψ�6A�L}�E�1|_+���[��8�K���g�A����F��/?�#1F���+���䮠<�֛��r���2���ЕV�������Z��[ow�u��Ŧ� �"b	A ;?ן,��sAY�+ڤ�lz�k����T��L��dq��z�����aD�P��M!50Kw���3�� �����1/`T� ]r��⾵��!���r+vk��-x�\n0ج�D���N�U9��J]/�� N���`W@q�;M6�*r3�1�����wk�)P��vmw3�^L+����oB���U�E����s4�x�n���U��v�����2R��J��_�ף�O��`�3|H=���۴+��$��v���^�`
��q7:,��b1X�����@��(:�Y�l���Ƨ\�[��T�� ��r]sB��<�#%�tay��w,FҤ����&�}��[�2����ؼj\����"��`r���/X��oԖ��� ���ZI1��t3�@��
�z��9 {$pzt<��+��åCoT�M;�s�|Ļ?����ŹD}���dFΤ��Ä��~��8�(�1J?���~���`�os�V�d��w�jR�VW��Î��6� iL�%X��}�̂|J���s���ɍ�n��(���F/P)�����C+W����-����ħ>wO4�n��'�dˇ��g����q3�'��-�s�a-�\�\5~:ڿ�q�t����u0/Q�� @���o���_��F>\�{?���b9.X4�hzd��NqHs4�mM`V��JL&A��dܱ�E��@��	!d��H�����^�#:�&%�]V=�A�5��mA��hMv�[^�S=ف���U��#�{g΍��CJ�ʣ���^I�Ս�\�aȕ���1�"]M�t�d�7�L���͘���<3��w�@$/��g���LϿ�gI�M{d�ٌ�4�/)U0k����Yn3!�G>� ~�ë���)��6Ўr� Tu�Y���'�V���3S�H��U'�sJ��p�L��Z]8K©b��E^�]bF��+XsU�n�EA@���O4P�*��߫'S�]������h��z�kYEz�W�y�E��d���1M���u<���-i�B���T����y�F���\�����k��<;���ϥ�"V��6ۑ퇳>���G������mu�$Ê�1�!�$qR������%�R0���i���t^bg�Z� �R�1��P�=)�À���D���)@�5T�[ⱕ	�	� ��(~Q��5�%SfI�;w֡wV�1�c3��VR81��?j?ֈ��C������u2p�4�����'�N!�|V��>��v$�<��m�\y�����%��A\K9��1��+G�Y����됆(�r��0�#�����-l��-��X,����!�M���	Ϲ��`([���p1Wws�-�Ju�����9)�C0u���h��W��r\{�m'y0�W2Qx��C�V��e��k�c�ϭ����8�b#��
��={ 
�4���_�$�aTr?	 ����q%�딸=�fD�
Ƈ!W���x��O+�w�]���Os��{"�# �?[���^-9�)��yZr�N �������moqS�]�Ak��/�֤���+��`�M�Z�7�'\.�'1p����m���#�rdamݹ`Oܺ���͗5�lҶ
	�xL���$���x&9s��\�=�}�j�j�֏j�\���^�B�A��G��'!�>�H���(ɏ�Vge���U���A�T������"ڝ����;�] �b𖃺�`����	��ZS���ǠZX�t;���|�$�*RO�k$��b�
��S�t�B9_1�ۿ����ڥV�'#���ʖ]E��f��L��6I�k�xV�#ғ��D
u���� �<��,|uru4�$��,��-�c_$��z<ga{D�,���|C�!҈��H�r-+�f��D���Y��b�Nj�Qkv4c�Q�s{ӈ���h���v��ў7@�0�'r���X�T��O�Ǵ���Q��QU$����q�O8S!��-}�����w`j��o#�v�T�o�����ۡ�a�TĦ
��:Z-��`�h���0�
�?շA�1/{��*�D��Y{^�����;P���C^�a8�a�k��W�aڷ
f��?��ů�0��H2�~3���'`S �E���^�&Ko�x���0��z��ֹMs)2%g����2��I��Z��<�����~�J���}y\����Ȓ9�%#�n�T߾��g:`�՝�=��+�WJfzXF�K�y � �`F��m��;ǒDJCcF!H5���|m��X�/N'�V�'kحs���hN�=�\�HBE��H���CۦO�@v��y�����+D0
~��v�f#���ci�n�I>L�鱒i)�]�Ǹ�fT6�>��\�U�#���l;��t���.�������h�@��ắfņ �O�ֲ7��k�����r���J����3��pI���9����_��ү���be/D钰8aI>TD�¹��P�D4��-̽ܽ��DL��ΏY@ ����)�p���}�(J�Ίi������5��~��rϊ�-��GC���(�H�>B�3�t�`H�]��P�u�?rp��O{߽`:�w7�c(
�CM,����|�û�Qhch�y��mv�BZ�ptg�,[��N,#�ƶ� �a9�l���'ӥ)d`'��Xe$�C�� 诊�u��A�9-��YsO�?0��?��~��f�H.��ö�h�^�Q�˒}���,&���2&���d�W�?�U�*�Q��N��6_�`׍�IĊ͍��zj��$%"PڴN
�J�i�SU�Ja�M^��B-��کsgķ����)h%�'��8%��CY/n�-�*��.�%wx��F*e(�`��1J�Ӹh D��5k�Zr�<ZL���8�4td0��}����6���T�o�� f�	[W��k[��	�#�aƚD۱0״ݮ1�`pU��@n#���aY��U$ܸ@G9��>�?��k+bl��R5Z�TU�2�Npl����@�%�<�)T_-^Rd��5<���K����[ 5�����w����:��-���|��շ���I+׷���ѽzqۑ}) �����ue�;<!ș���\^�n���N��Y��&�Z�ѝ^���=�@��AX7`Qq�n=i�,�D��G3�/8�'��HzW��ZV����~�kd�F�y�g&�C�	҆�<�?6�F���е�]y�����r��v�����M�&�1��_�`�-��^�*����O7k����1Z/���6���{���m��N�kj�x�s��+�1$�<��n,Y�$���I�<o?�D��"),%���T7ڭ�V袛�m�p�c�_7�j�R��!D��j���'R`w�!bV��2P?�{L*�>.��m�с�m��#�Yp�h�0�q���t��)dڹpZ��&�]��� %����n�ҷ#h[W�K� w@ǁwdwۭ�>}P	�O�>@XY(�	=���l��(�Cg�?� NN�ke�9:Qm�d������[�2�t7��x���9  ��`�XF6�m�?��-B�����W��c��j�8e.������C�6=VRWi�|��̼w:a2�0�lȜ��u�b%�3��.�8�&�3(�vjJ2����q�_� q|/�/Z-Y�n��A���̺��Z�.PP��)`�'��Iƭ�o��k��k[�ަ�(O�O��0S��k,��qzu������0%�NFl��~�e������M]��1��L��C�ث'Z��Hg��[��=��G�f#�_gE�S��H�S ���n-g-��ۍ�բY�0��$��i9�:�m���e6k�Y����z�tY�P�n��cf�2�f���f� ��D�|�d�7�M��p)���%�B�횽&#/;ٟw0X������W�&c�|�?Q�Љ�8j�G�����+��^VW���~�2\|�#�ţ�z.)�����ƣ���m�92���γ�Wz�b�·��V�U*�1�{
9��j�H#�X��G���3s����\w�h�vS��m�v ��?�u1aumr��̣��&�Ш]����^���)m������U&L���������-@L�b��d���oc��1&�#*!g�{�(�1}��W�+}�an#��Yu�т@�ԣ��K/�a���*e_�M�E��ع����kzwX�6wT{�#Zd�C��rC9�V����^cx0"Q�õ��~�"��2�n#�e�l�\�?�^N�9?�~9��H�0�� ��I�����1�.ex�>G2�;��;�d��v1ܧ��a}�9����E��>���$�Fͻ*v�� �p�nT�8��z~n��Q˲&mHִe�\������Sv��W�K,���z�=� |L����J������
��Y2�;����/q��zҐ��mg�Gas�nY��L����l�S��p
$��tcS~� |��0^�o��'�cƲ7iK7�PO쿅<Ҡ)t6�����L�-�C��d0![ǜ�e�J=���?+;��9��l!�*s�Wcb��[�R[�#�����t������0Z�6|�&�Q�"l�����h�� W����K��iIg{���pø���p^[�h�+кT�Dx�M��XlxVHYEB    4f27     d40�?0���7�/7~�מ�ظ����E�9%���W�c�����oG�?q����O^����Le�]�l��zՓ��m�v�G���W㢙jM�S��5�BZ�����I"j��F��7�,ؙ"�f�D�ѥ�ukHG�Q�S��)~�d�bT =A]:�K~TKIfu.�?ϔJ�a��vX�|��G���w��;�]'Ǹ៪�%�I����<�(�82�g4Y�	cf	��c&j�z�r��d�51@`�ɷ�=(�������#'!fb`ľ&�@)�[v��Du:�_ɵ�*`��*��Nu5�6-7�� ��9o��!�!z���
.�A	�āAo�}��[a�LX�"���V� f��ܞ��8�%��5#4D���Lk�T�{���,�d�y]����(5D�x��9�� o��l�e���=2���&l��g)���X4��x����9�YNos�	��;��/����OB��(�A�/Rq�v��PBV�&����M���;���f<���s�Բ1nFv��%� �XAf�+�"T��d�ī�{/˔���I~���B�ek7��7�锔�nNQ� ]���b9Er��<|���e��b
Α�\OT����嘃�#��j��ע%�#[��J�7�y��3����mC4G�����S��>�����43�Y6�>�+m�b?E���@��3&+xh�вc�����(E�	�: �R������>���K�>p_㎗Bz8'^^����2`����Qb"x��5�P���"gz��Z�#u,�αǏCs�0�.�-��@e�ا���ǩ�at0F��q���P7����X2acc��*��Jr���
�K���M�'L#�8�[/�!̓Te�KO��5�<~�!~��2td��1���Tq3ɜ� rf��g=�%H�j��1i��<�t��I�>Z���$�{�7�e�-�yRS�����J�1�.��@��m���Bv]�'76�th��P�����(����
��-��C~�Z�A!Dv��T�~�ۈe�$��<}���Ðc�ET�m3r�z���M�4�$�f#A���ND���U�ǇG[2������J���}�c#��$�sf�h	=��t�K���ޚ�e��u��<��:PL6��n^���2P#7v�`���_QF��d��p=�����^�1=�5�iD�0�$���T��рdxA��C��N��i\�?����xZ�hg��wۃ`"�Vv�jpb�476S�.24廈���q�{g�1�JG�Ѧ$�V6|	]H�RZs�=�(<n�;.��rѶ�q/�2��V�c��i6n؛��X������=��'	�1��6��XK�:lN��(]y+�8�Eȑ3���> J�������:w�nH�ƙO!C��� &MIR� �[(���a=}/+��ڼ��E<e�i�����xaF�>�ҷ`��L��~�V5����_V�5���"z�}���-,'$�f��S��I?r�Ô�?��/}/����B�%��h0�o>�J��7�������r~�P�m��N�G[���R����`�C��ر���^R�C��g�M��k�	'<>X��"a:�]����x�mt���W�
��-6g�EC��>�t�x�/+�G�
˗��!����	�\��䧱bE��;�Yv��R��Z9ԏs�L���x	:@Otp�������0���A�ch�3|���p	�d�Q�џR�n*���9w��R��۫`myIl�J��|����'M�X�ͺ(���k������ F��p�QD3�r��n�6ٲh��#q	y�]��<Oz%�W餻ևB�q����6J+�2�'���*d~X�2��n��XjL��b�_�o�݈OyE�����"�_��p�+�$�'���FE�R7D�J��[�)6J�����Y��I����l�ƺ���(�]��P����cx�`��zO(���U&�7���	�+n.p�ݱ}G���½���U+��t",�۴؅�=���O�T�-��z�9!���K�f[Ī`_T�0'�T����&�/W�	bֿO�����P:��Η�Re�-D\bHs�Ժ�h�kNQ�*�F"�a����.q�y%<9���Y�D���9F��##��gh�y����C*�bn��d'~�ۤN4fmt�HC�\߮S� ��+�]������^kGhA��Ϩ1A~#.b�~�*��Z�w	����Ԓ٦a�=�5W��|�g���FP����.�Ąx�flɠ��!��:8���Հ��}E�1{���[�|�x,�:S2L�@xKG^nւ���I@>F虶��rzV$�+[h��ε{,e��	�<��?\Aj�������_�D���H���c�;/,�|�3�1aeQݿ%,4$DVI��w��#cq�*�ĠB��6���C��dL��ƹ��0��k#'Pk�47Z#�nxrk0���C�|��=�4;9j�	��5[�&��z��@��'�9z���n�s	���N��@Q~8�$�-۾�����x})5���]�� _�;u�*���h�51�����K�L����A�9�����z����-��MMk�=�(y}�O5���6�O8)f9v�t'@:mڔ!g=��V�K�s�3^��Fz���t������c3A:�c�\e>�l�Ř^E�8��� m˸�,�)��b���)tAv �T�fK9#}�����0��D99Й�]�{�w�Tqo�<>���EW�+w|$�\��s���j7&f�{��r�0���F28���t��7��]�� �H����ͩY7�P�&�~e������(��z���� ���7v �E�po�����RĀo�m3r%%y^��$��~�w�u2��� ��`J��]s���"8�#V�. 7>�o���߫�R���X�]W�|1�Bt�ɳ�����R/T˱Y��	r{����e��-���Z(����X�%X]FG���)�c~ϐ�~�[��/\����5�O�bϜ����Y�:[h���{��=.�h�����nb�B>��2�`�o��I�|j�4*��E�	,zi���Ě&h�E� ��̴sP�zuj0۪����Oq ��
��Լ��|;��[�B��]�sb��P�
|Sn�y[�Cq9���u�������r�N^ah$�m��Ol���o��0�[%uV�E�GaF���L껮 ��ؽ��a� ��6����a�TNF����:�i�3��q�5�{��C�D����l�RP�H��m^Z]�M)W�%���a�y��2���Zq�1���X�|�>��\�|x�nf˂�!s���	��EA��]��