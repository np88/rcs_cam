XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��eZ��E��M_�"�gԗXx��y/�1�%U*+�C���,�̵F�ǵdbĝ�ԡ��͇�}@���D���V����~̕��.�+i_e͙��jŞ���c
�4����G�����*#q�WM��.޴��$�5��LK�R��
�nH1ܺۘ7��)n1M�I���@���?P��'���x��%�����R|�JUwx�WD���k]�nt�LU��p�(z$�r8;���Z�i����u'��M䜿(��8�@�#�H�����T)/d����`�@e���ƼAw���	=��k+�{���mW��Jk�R`JU�.1����>3@����0�O\�:�)7��tT�]��@������U\�!����]S�VQ���<X Ћ{�D���;���S�¶
뤶�7�zox�K��WI�fw����$���Ƨ�h�='�۸�p���`+�âu��u����L؛��ge:�F��c/��}A?,-?�<u��;6�U�9.�8��`D���}�]B+�ɭe]I�Em����d�LGP�?�����qN����L*2���I+i�%�i��g�i�)ʆ*�&雰�"~����hm:\U�z�j�Q0^��� �|��pC@������UB�Kp��T@�^��_��c�>��0���S/�k [�8�]v�j.�h��s�\�%��ؔčC���Y1���s2�A-;p=�=z�/�$P��"m�̹�������v�9��!�eXlxVHYEB    2533     b00F� ��zG�<���e�9_�Ð�AA媐c�����f�R�ㅦ����vYE��J�ǚH�^qr�|��H.����"t���~K3��CG-��B$Ai�s��t��=D��!���]��
�E,W�y�v���L0���+'����,��M�Ms��s*I�fE�h���\H���?+v�Se�!�����Y��)����4��k���PIk�{�q:r(|?p��w���x�������Q���8� �g�U�
c&���2�m�[G^j7H�Q����Zn*᝺�j=x$�I��GX_�o����a���*6�%�|E��ǚe�=��@�T�1�AY`S��>BF���vW���v��'���ڥ��iz5�=�1ʡ��z�>�̼J(�F�3�9@(���K6kV��sF��1C>�UG`��=B�|-ъ�8.Ø�e�c���^���NC�\�G��c?����������2�X�gy�bq�v*���e�v.�3�L��Bn�ք�����-�zhw��:���yx���"��=Y��N����/� �O@��P&9�i�+�3v��U^2�z�4�>B�ۼ��ǢR�#W(�o��<=~�N7��?��,RQ�������jO����%�mңF�h�gV"���5�a��ՁB��FFM����3N;���*R������b�x?�vwu��&���.U��˝o6��~���{Sjm�>�Y�d��7*��!�*o-(����!�}��R>2�Ǯ�5��r�a`��k���t|��ve������s�kf�vg?߈��G%z��y�4��"� +2=�ˮR��}Y�}��Ŝ����>6�C�_�/��'�U�,��79�;k��Uh�↸��6��1jv��!�z h��V�3�W���JW*2��C3(,�,R�0ҷ���:�� MB��$J95w"y�` R���
�x��bm��Ӫ	��ի��L;�z��޼�2�6���0LL����P>�@Mt��G�ݿ�ੴ��.@��x$GI�C�9�֜�	޿��m������M�:g���+���!�'0CA-.��ᷳLQeU���\�qݎ��բ�#~�W�i�Ff�����[��NM���2:��O�jφ2�\�:to�e�鍌������F�:�ՙW�1-WW�h������V����D��{f�x��W�6��n��T��/=ȏ�-P%�ţu�V�`O�JH�W!ޟ��W,��m<�x�s�����A�r,p�`и��VP�jx�Ș�ɒZ\�Z��	%ĸ���"�9��j$}�B�I��Yb*x����!Iأ����&X����	�}�	�Y~0a�7H6�4��@���]�#6$�3���C�3���9�&o:f� Mn��H&?Qp�{p�� �X�(	GN��.]�H��XO�@R��[���>�yL�n�PγmOj��Y�uKˑ�тj��نQ['X&�HA��3^�0�X[G�Uɝ�&�h#˲�n�lRr��7��3Yn~�/c��=�3Q�%Z������3S�b��X����^��L�P����F~¶d8��0�bg�5FC�b��t�!�#��4��%���>o�Oa24���l��Na�6�����Bo�!6�C�F��x 50�3��%�)q{���V���oSf���F�L7�ܯ~�bc�m�g����.h	B��	|��6#-�x��NJbsP�gL��_tR����W?;�=��t��FL=̯� �l|����+��+*c�មc}W`�܅�������Bd�JS�br�?�\�&1 χ}Q�����M}A�����`uZu_�U	-ã�ü�uhK�HNjYrf&L�R�%y�?�����Sa��%�d9b	��D��;%�j���:����P�u�t����V��_{����7�%u�s:/e�7�壐�)@���G���2 ����L�l�v��[T��7Տ3e-_P��r#a��-v�[���������M!{����B����u��~F:��̣���M�/z��V���7a�y#ɍ���?O�43�j��p��HH��aح���8l�F�cQ�cE��q����U���s{�ƛ���X��о�R�/+��C��FUU'��!.��2��ݕ+rB2!��M�n6d�����e�azKu�� Q*�k����0����Z]�V�?�?T��)���e!V@���� �o���/G)��J�jk�MF�� E�sp��},{�B��c��2Az�����O�_R�2�F�N��\�a?��F5��$`�!�f����[u���	�LhQ�B�r)����e�n� ��);'	��!��g�ǰ���؅&D�N�}$��w�&��1�0%�2�Ws`J�QlFV3���Ipm�&�1Q׎6j�Te�������=���w�SE��dw ��XZ����^�]�G�`��vn�
�e񑷧� \�`x�1$��*�-{�>��3.V�x@?�߸����=Zʃ��s�_>:O�u��Xň�ߠ�����9�k��1��g�5�{fa3��W���?Hyr��fco�Jn��I�y�����gI4'��,�gRoE�
�7#d�6�`w���Ϟ��;f�$l���^5�d�����p0b,S���o<j�l6�q-��{���Ը����$E�a@[eN)�:�^�N�D� �d�]�Pl�-����)A������w�IK<��4e2 V�w�&�H���CV��1�3�1� 2m� /�:���B
����i���