XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Zˣ~^�}�ٲ��ٖ��b�C(0X䡪�H���޹�1�� pe�u�A9n�6�.��o���8�Wm��6H_�kN��x*!T.���(e~G�0R�!��Cw�y}yWg�Ck��8�{O���7<Y.
H;ya���/,�Oǵ��7�-Na���ҩ��I���f�7q��<	��i�7����d�8:.��\5�H7��*��<�:���ʗYשb?AH��!��N�C��pb�Q�y��!j��� ��Zj�r�<�:�R� h,:�nn"���N;������*o,��!b��{j�;;5��M����= �5�+m/��կ�'�B%�� a �8��
zq��>E�$��wpv�3�FQ�5���cۣi*��2%w�����)�sz���Ѐ�@�l��9�V� 5	
~-r&����Q��k��Z�����'@��	�z ��]�c�D�޺���W���8��w�:s��_v�Y��
i�iW��ع�|;�X��d�˶�i�e9YH�k�<�oޡЯx �huw4� ��жE{\�<��?1^:�AzC��{r�/�����E%+	D�r�)$_P7��gǲ؋A�=ab��UV�F"VCsf������o���~��͎2|���K�qXX ��$�=b��$���W��A�}!5�y"c�L�+��qԭ4f<�	�Ke��} 3c�3Ͻ�'4'�&oS�"�Z��B�Yo?{�����Q��.Y�P
�>ZRO�<��`3nKo̥��2~XlxVHYEB    fa00    2d70&�������'�
��+x�|�:m��m��b���\2���z���{��:n�s#����=��#� <���K,E
�/�N���Q/���LD1>�+�qz�WO���g���7��5��iٲd0���Q��Ip��^��	/��ECMP��}9���@`@��笴d�4]ƣ���2��4�{}��;��	�]5M�4��%4,��]���9f�3YlP��j��ԬV��ەH��&��l�)Q���D�$��_Mj�
�����u2�43�B��]��4�H'g�, ���j<�Xye�/.j����I��3$�E�������h�"A�<�nW{�h.L�J��p�'���O7U:k�y ��5���g����ܵA�곗��G,Ȣ"���������F�N{���O�A'�KV�����o�VDj���s ���bG���Pӭ��i���
�Z�|S1����(��x$A���XjO�[��=?M����eؕ�����s�TN�N� QV�<Zq=Ѯ^��3���[�+��Ĉ3�$-��
Zs�-w���.��ܲ�N̓�����g1��O�|{[r5���cb�+	�}?Vŋ�B��1q�FÈ��[]g#�U�¸����kЈ߷׍�(�m ��M��c�r��1�d�]�-%xn�c8��#q�񫋖C�V�}���m�4V�U�'���<��0S��%?P���[����xjfD@������?brеD~�L����>�b�� >ϴt�jq��h�ԇ�d�+K��C7ƿ��]��yt[C��࣠d�÷.�(�|�z����Z?a��Ce�����c��z�v��M�z"k@,������g(=��Ԇ��g�T����n���&���]��r�z��RӠ�iv�R<������*�H[k����)�PZ�Y�l>�	uY�]0V�����{םLX`]z���ړOW�Ի�D\Z0Oː}��V
K ����,��8��+3��{F�+Y	�!�U���EZ6�RbV@}�b&��u��ɰ�A����!{��yk"`����gZ
'
O�Y{����H�S���JO27H4|��~n�˸�\���%�kӍ�v�Q����.h���4�`�y/_�R�٠��� ��Pӯ~DG��~{���)o�g��k�h8+�����z�b��U���'+�
)���6G4����=we�1�F�>pg�7ju�j���Vƴ���(r��D�C6w��LP��񽳭c�~M49SM�� ��t`$04qZ�x\�+ax	���[��7ma�e���1<ɾ� u��poQ�n5�b��4�zm�#�>����n��p� ������j�I��
*i�Z�<�9{�J{H�����D5m���O��Vd��\�٘"�d���җ	h����9?��z?d���>_�>F8ɜŀ��qUeQ����+"�`�bC����G�0^�J��_�8av��Z>�N�d&|�$$�s���4
�nFpg{�e��7O֛��u&$U��T�J*��x�����3����k�#�D��`��l£ԙp�1pM2x�y1�1���R��ʡ~��z��i�*;��3Ҋ3��V�)�|]�
�[G�?f:�?�ݸ��Md�_�Ok�Y;��Aa
N���u���m��
U
H*h}�04�]he�߅��p�R���_,g7��S��S�㞷��C��`�J�=��Dz�"���~�f�.���˫���x*�;�jϜ,U(D��c�����TP�[]֤��Ґ��a��9�c�V��e&��o�F$t��?�j�u�"G��R����pV�X�ߋ����ݠ�z�T��f<��{�=��	�^�\���-9����'}�c&��E-<��$����5���5�����������XmJGɸ�'�lwpC�Zv�.P���w42��[�cp��7��9��"�1`��{���n�e����ڊ�'��H�F��������21h�c��赥k2���J��c><6�c�T���#>�F1A:5�U����~g�
�l�Ϣ����q�R B~��Zb�A���y� ����֚h�Sa�-/��0p♆dB�<��̶W�N��nH��WK@N+����~�-�5R�ޯ�'��= �.g��cMé�;���
�q�rXH_�/6�i�]��|_�m޾��bQ��졻D��O()�}4ͨ�!�vX6���-���ɀ$t�=I����ێB�E�Y�������,�7j�uJK��
䅌� ��%��0DS�Kc99��-q��?��R��uB�]`s��B�i��x�;���,���tC�����1����i̷�h)w��K��6�8�;wi?cd�,V�P�>��_w��R��姶��G�?um��l�6K���f���-ZOM�D	��<�?z�~�A�W@V�9h�bG+)��'TɷG�Ki+Us�����K�j���է�:Yx�e��~�ٽT5�C$l����+��9,#�� @�+P�l�H�	�ܚ��؈v��~�M9=0˜}E3]%P��&�S~֨�J�*̐g%k;J����;e�\�t���:��}��1J�ߥ�%���8u�Z��;$�� j��!��#yJӶ�����;mkV%Ќd�#8����@a�<��MqQ����ɯ@1��l�t�>��7y���E����-g�up|M��������'�|��k1BaڱJ�s���_l|�U��ϞR�`*?�2�*���!�y�Z���@RB���W�d$�*�ۣz�r�ڐ5��q�;��V����zӈg��}�z���D��g�˒��u��>M���(©��A���B���~�DZL���0�li���Aߣ&%O�Lw�a�PmC���;��
�����_{!TkZ|i"����S5��w��).���Tx@f��׵���U��z�s��z1�ߔ.�����WHB.G(9i?/Ϳ~�e�R��4�X0\�㪫�F91�N��&����OɃx�@��L:��f	j^����Ь?�������N٫��k�V��Sf�9~�0N��0k�%�P��o&��c,G�W���s�o	��]Ω�
Z���l��FէAWyeO5��ͧ Ҩ���R�����p*m����s䨛�����"re[^�_�`#�.������"�
��>��On�;>��IV�	���6����m���`�t�����n�/���E�t�^�Ϧ�O$���4x{k�Ep��A'@mF �&f���ri�m}�{�)��ITp���_w�W��ٮS4��?��&9��S@9k*�uٛ�&HU� !)"�֘<2u�M�����3i�SC�=���3;y�s�+���>�9 �︅AK�M[�����(N��|�.Pz&�xf&ʭ$���s0W g��E�+˴��2��'c�i�_r#
 ��)���Bx��zh�u�}P/��m��e�j{q�V�"�wWiO�X�G�� �k��T4���ϱie�������r�qC�E�]�]K)?}#��cd��[��Y)�/f�Rʼ:���%�;����S	�!2�_����a�P^�D�Y O��.}w��2�&����
]a�&n	Ļ��2�,cjŇ������"�E2i�����3�z���jк�q7�faRt����N]l���^��R��/@���T�O@���|ߊ�N[�����ѣ
w�����]�{�w�����_c��I��o����;ő:Ǟ~���;4|]-����6E��^|��uE�s�����7����ug�3FV)��w^��8�F��gi�e:%�1<�E����[��9��T��4�KV!�n�S�������O�,����G�L<��5�ϐ9�N��s��K� ?v�c���Q��B5z`�L j-��	��F�}-{@2C��H��g�6B���.���J7pL2�{�o��͡ΐŉWѓ�1��2�(�}e�6D�?��-�U���X|HkC�
);��3���M	9��@����N�0��g�Qe�L� �����8�n����c��P��fhwT��6U~X�>.�%Oo�3V����{��Ѷ=�J�CNl��Cm��Oq+[���R�PѾr�zC�t�q#=��f�)RwV�3ֻ��3�x���t}�=�ჲb�`2�5Z �P�=�6�4ۃT\��gCm�c���g�B�#U�U-3�9_���uMJ%TH>�8>���q\�Ŧh�����S��綵3�-�+'w%nfI�A��NZ�(���dY���ς`�|	ި����Y7m#X3H҅�j��fM[�O0#�6��YV�-��mK�r4ԏr Nqa �(Y!�gb.]�M�
O�W0_����|�� l���+�M2���}~��'�34=��ۻ+�:Y��Ƚ�K����Ր�n=;G��S�E��+u��Q�����7���pX�C%�4���h�[ܒT��+�23����)��k�]�_��;�MJ���PӁ�w��A�����X��ā�9�2�!�l�=�8�6��e/Ӹ^G��JG�pb?2���	;/yW���4p��x�xʹ�|_�����9�vX��j���q�^T�h,d�k&狪��\Z�%�_@������3#�E��P�EX��=�ׯ��G��nB�:PT3���>��mN�iM�������y���`�4�I5;���M��-$n|�1.~jⵍt �Nȏ*�z����N��D��T�.��͘�!v`�xq���v�9|1�N�3�f�i+GE@����*p�mȯ��\JY�K-b��tX��ű��z��p�w�8����7��2R����S����C�Z��"��a2_��*�&�9�����y�HD�I���3V;*�*���?��S�(��;/Y��XGr��x��T�\�+���Nѧ���k�%�X��'��inA�rZ@�1P���5�A734�d2�%=��c
heBԙ�F����Y�0�e�긒vgzL�q���Ԋ�����S,�5�g=j ��,.��s�2{�|�v{�kp��j2�!�.�a@"��@�����Y5�s��`�H��GG�����^�<	��} ������:�����_�L���w����&+V/���BEֱ+]�E�e����vC�g��n>K$]�o�n�D~���W�Q��ָ]���`?>'2��^Y��c]m�ɳjZ
J�����*x�(R��*�Z�SO԰22�gP�w��%-���.OԬ�c��q��`��lh˧����70sk�u�^��|NWc������R2~��hE;�ܮ����iz[���	<)y�Ι���.{G�9�=ϗ��4����U�m����؂�"
��]��iW�juq�g����꘽͇�}2���W��S�n�+���}��
�����3�5'���"}�,0!�̄�4��c���ǡ*l��Bͨ*̫����vI�zƸ���_�8�U�C®8Jo���z�q���Br^�gF�~^���C���#�������f�����V��[�.bt����(��Y�#E{\<((wF��3�Ֆ�ߌ�0(�v7��&�)��)tūco���`�P;j��^�o�0����0Ah��
�@�:x�^�5[�E�}l@e�,~ht�%]�"-.�/7�eѰ�!���A_��5Hh9���k�WmN�����Zn���J��\����$��<'fn�Ӫ羉�z�e0��k_���z�A�ڟ5�4��S�z�$J��T�@`���>0��#�;��,1��p�� k)C^��F>��n��e6/Ͱ;��:U�g��:0Z��ʎIo@g���W˞=l��-�=�n�l���
�[�c@-��#��0c�V7�)�+����k|��Sm�b�󠀛�Q���%�=����X<�����^g����qa����㓬��D�f�������]��jG�۷=z�Oz�0�A�J;�>�d�/�ڜ�E��G(�c.V��-��1��*�M��u�/�y"h \���*֫�+�{2�#�B\��$658Uh�r��rV��_@�xSU㪕�@?#q�� �ԓ�/��o�{���3I�i/i����
W�y:������=0�?2 ����1��=�JD> hHi�ݽa���PZ���7�=�k���>���@]���샣s&~X�׫]A֋}�C���)��[�c�X�~dr�\ٹF���!��7I �����8��;,>٥8.��1��MLQ*�y��v���}uH���ķ���
[iP��v�wӸY)]�솞唥@��U����r ���ӭ �/�=��C�Z��5��t79��s֪D���k��i0L�.�Lp.���
�]	-�1�[c���Q�L�9y6���\������e��>�aRl���,�|R���:�3���i��j���W<%\��ӂ#)r�[�ݞ�H�Zh��ز��֞='�=�W9�mjJ,��9�U���#wg�gKLԭ/���5}�}��u��k#`�"�����D�)CYo�Յ������W��6w��q�fp�߫\�C������E\+r�sh��bҗ;u!s'�2^�}���u�]S�4�`%>�z�hܬ��-�#�`���c�ze����?d��	c.���MſC������ ����p_`�{�v� N�&p�W:����\;��e������"S���L�Lv.��$f�SUIG1�*��Ӱ�ɹ�2k��w1�n�5Y+a����M�r�:Hk~�*��Xj�n���N���D^�429?���K^C���R���|,�Z�������T�l�����U���[�X�6}�I�j����;)�Bk����I�C��4��-�}10kP��_+�al�;L� �/��{ �T|�w�^@��������o��M�J
Xr� 2��l%�������?��J���W�y����`V6<�g^�����f	I�'o�FHY'_���C�՝$~��a�f����L�����v���Z�n0t�$RG5������2D���ړ'Lʽ>�Z������G��YMM¾�/���U>�Y���L�dU{f�$��83�A�[uQ���Rڎ	����8����x�oሽ���0@Oc'��j�L��1������MʺG�z����m׫����`������
7R{l*l>K��0�/%�]��d�l�j�k[v�Om�� Ɔ,���F�SM7��fʫ_�"���	��!����~ͧk㥐��4���hZi�$heZB�ynT���Q��q	�/�q��D��ޞ�ٮF6����zh��.9f>�J����s�/K�Y�b�j����^�)s�Wr�Np�0,D���'���K�S��B������8�[�K(ev�,(4ĉ���a����4Բ(F�� ���^��8aC�}SK�sF+���	� �x�����&�`���H܃�0F[���t�Wq] ���������nWD�:$�K[֪�j����A�����ن�<����@����C3V�j��8�c��ex0,��#$�����tW������L�xF��D�_� ���[A gWޕ�8��*V��zD�Ã�}����xd��4*�ưsWLoB�Ɓo{�EG0XUlgyw���e^�%�2�I��Ç��h܍�Q��h_�D��9__�Ju�{�����s����f+���VG��jŀJ;�3��13�������E�����RA+ftw�2F�օq���!:�����>a�RĻ˯�/��r�+c��9c���]��K�~��n�n���崰gU��&4����y�۸Yv�xD-�/�,�Z	���6w�?�l��N�"[�*#'d���r�_Q��ox��\0A9����ޯ����I��3U��cQ����E{�ߢ L��K�K	�٘Qg��)��D��� �F�a��EOv�\�#݉O���P��n8c���?iXfi�,�d�7�--31�c�4��"\�7\���.}Ԛ�!�wM�������
Z�RM���'z��l�� ����M��G/�iT���%c�GX�i����}�ģ���0�޲!7~X��Gx���������t.�) .�(�@}����C7�%�	y!N񻙝n�ѝ=I�gb �bz�Ú�[-J�q��*���;)�5�����Ρ::��d	U��A����Ҭ��T�r5^?��%�R4e�<QХ��?O��C� ��w�%���Q��-��>,�t�<I18�|�R�X�I����{,4'Z�A�A����**���*k�ڀP0+/|H/�K@j�q��ቛ��e�Z��@��G�9�)��lh=�d�ВXZ�Wzw�9B�̨�ib5�uZ�B�ٮ�J���#�5�X���+�������@c<@U�I&>����v��Ц�)2�Ʋ���xw��B��$"J��(�u�8�|�!x��{��S� ��������,E �}=�<��
?Lp�a�� �4�t��"���Ң�&.�*��W����,�_p	t��c#�&�6��n�o�=S���n���l�������BHg0Nv�e�(��ձf�&��C�3 4��/v�?�"`��Lc��L�5d(�0��cx���o��Ks�����N��r��`I��=���h����?1�g��
��3�� 	K��j��.1M��ȭ#o��A���!�^!�ɑ��r)��5���[@�"�G�ر��PQ �V:���V�|S_f���!�U�{�k�"H���]a�!Y�����(I�����bMES��66��5��V&+�SV���'�D������S�zQ�Y���f�n3ܨ.��%���{�y�U���o����A�d�K-�#f�KG?R��=���I��綃A���� 7��k���݁��v�W��ē��̂�ܰ�p���D6��٠_=Z
@=�_��a��3���
�W�6l~ȟ6�	��p��D	T���5��z�4:��o�@��
�5o\4K���r\V7�J�6�RYp�C4q�SO�o����G#`�}vD�;���rq7��:cl�2@�.
,!S\�q<��@��A���qA�w%Vc���k�]b��n I:E�z����L>�ɰ��>s������)]��ϪM�e��b�1S+��e���ъtek�2�Z���xJ���h���/rR�T�$�Oi�9Z)a���MQap9c���n���2�@
��{\��qFW�b�|a�ٌs�iؼ��Y�A��<�$5�Ӆ4����w^I�~l)r�X��(�R P�yzcs��64}H�._���9#�0��a��K0uy�c�h�
���JU��y��߻�/���&#�&�[�=�j3$(��nh)-�x� ��L.��̧`��NG[��/�[�,X-1��ftӺ��*͑�1�]���`�cC��U��iL�8�j�?P�8��fDG���-�w�A/ʗ1���	���~�SXo��}08�WZ[��`���Lh�_NX�Ӄ�D& )�:�q�2tDinxl���?�)>��­,���ύ����&�|#�uX@�?9nŋ��\4�~�:P��ɛo�����=J�EG��_WN��H���I���d\f%�L8�pS�4��[�x�]��^+Js�z�l6������� ��bULb�M�I7i���?�ğx�#�v�*@\�?�����4 7h��t�l��:�S�n��R����ޔ+���`E�c���0M_�3�N�Թ-Տ$�BLs��s��*�$]EZc�}��0������GׅZ��ʪۮ9a��+
��6�aA PQm�>�O�o�?��� �>����d�<�c�&:uE~]�6��ʗ��T�����8%v������W�'���}�m��MI��CW�x�,��0;�`I��ظ���yB��m�<u����Z�"���T/�Y�MS١�������*�~��OB-���)��2<�4�����B^G�$ϭi��� �O)!f>���f��B���r�a_�z �5�>u2��ٲ�
���}nA�����t*����pFS�ŁL1�a�r�\�<�i��0�O>󉈜g�İQ�d�j�[�w���~�Z��#���k��� ����.���uDĔ�x��0L�B��ޜ�ŤE��co,"�GKJ��|i[���Zz:�`���J��<�M�{���D�g.`��K���tP�k���[��:��>� V+|��>�� R�u �A�Q9Ӵ��_�_��T�����T��_t�`����SP8�% |1�k�e2� �c�2�׊�HQ3�<��Q73`�3��U��{�7����D-%Ĵ�З�$�w�X�Y���/�+V�u��
E,���CRޔH�|#���7JEs-L���k58{bno3߫W�M��_�<�~�]�urs8�bԸJ���T���\ac�z�	���W�kC8;l�qG���66�����P7E��N��b�n\���'1�E��+䞫N� ̷j���aa�q�Y@�(�A�g	f��Rk�q���o��a�U7���rr��sڪ�x��Rbq�ɞ)�-Hi��z����4 9����!ֵEs�(�%N>辏	��
vf�G����>�T��}�T��s	C��J�bu�G�V�(��@�,��BU�����톳v���+��!fS]�N�6|#7ҼӄW-6�s+bId�LyĲ�Lb�#}��VU�k9n��+�V��p��U2^J��-W�/�G�N4�/Yu�vhd��D�6��k(ow�SɾqRO�'�d���?Z��S��7��R��́����H��庭�7��u��1i�@�=rڕ��;��g�-Z�MaӲ�C����b�>��&��i`,l単t>��v�o�0��O*׺����߹Y�QK_�z8*����,Qհ���ն�W������+� �Ԛd�o��Å�����	T�+�M"N/w(�?�(���q棣��^���=- ;�)��cƏ��6|�lH�aٗP��?(ǡ69�~Q��_�s;E�Ka�3�0�:��`�N�
y�ò
oE����7��nujZO��c{��3��v�A:��̶e�k-T������a�5��|33�^u���t��`;�K:�醸4P�B���	�����ܲ�^zoID��g��M ^(��㢓r�=�v,�-�) �D��N�/��P�g%���H�u$���刽��L�{�t\��h��C<�����p0h�����R]����_N�)�'��K?�_��R5Cy��c{h�n��;��z`w���s�]��e.�����o�>Z��آ;",x��̀����tMUbo�=���+y�_J	ST*�x�3͇"e�%N�8���+g�F�C���/��aYqeU�B��g�(�Q�f~���Ƕ��q�8=�i&�?/���~� K�G��+��=���'0�1����_ϖ%�vP2���0)����B���X��߻���H;r���x5XlxVHYEB    590c     f20�}���uL�?�P�J���#���.sr��5Y��*�~���5�E��쀰p���a�6�+��g"� �\>	E����^�e�*X�,q� EVCG[S��ߪ+�H�=�B?k bo�"9V�)��m�V.k���錘�)�����6�o�jŪ؍�$���x����<���V���3��C�"�d)t�M��92^�I�xR\���:
#G�L��K+�JOuE�y��< ]�IM���2��"q�ky�o�u� R)͆�t��?� ���mRw�4�y���W�a�ѽ�m	�U�F�HH# �A��M�X]j1�&���U��}�fN�����ئ��c���x��<'�oT����^�a�Z(��xlc�4�s ��4���Z,F�R���[��� }�(�ŕ���&�`Q��[�1+�V���Ǖ���j��;�B�:s��?'��Z���lC+Į|�<��ȹ�Rz���J���T0���i����=g��[*�ER���*�ϼs��b�l��7�?~�-ng`�A�?���V;RiG\�u��"�Q��p��c�"2���zF�DZ�*����~���W@�3{BYQ�j7C �g3�����K����Z����#����e��{���N���Âm�s
�P�+.��>�eCYŻ�-��+�FlU���idDRߖ��ƞZ!α���4��_��qW��\�pqe2H���	����K��q,
��sT���b�[��z��}�^,ݺc�B� V/�i3Ry؋� �~��h���:�����vY��.Am>�a�ݷ��f�j�]Y-p��w�®=V���Ou��j�F �{�a�uoN��\e�����]��4���3M��J㎳J�Up��4N�q47/	9�U�3��k.!�!�B��6E�ĥ�X�{N�r��u��h�oI��sgEw['#�XS,S�C�ʡ|�J�5=ʟU!��cݰ�����=$PF��a��t�ߌC��R�˸�$�_��vS�c��½�6ڔ�~�s=g�-�Ӱ=^	��ET�G� -� ��GaX���(6�(O�5*�U��n��-�E#QR�@jgJ#� ̩�j�٤�����*������� ��� ���V�W6��7�xq�6���D5P��8��U�7��_�0�R_1"�zqX}�֪%)^b��H����:����꬞�w�����)�S���r� E�i���4V��LiRk�r'X�I�x-�f5��{�����v�<R����,��Ոk
Y��2�.�q�2�s;�$�s�} >��w�O�u�ؾMߎ I�s^��i/wL=��AkD�oU��C�9��n�~^�&͓N��;y�ɧ+��!������O��L�W��b�~�L`5�?���m�կ�����Ѽ[j�AI��<�{&�~%'������h��I͝����]�0��R��T�	��ɤ_]�~�j��|pRn��	�T���]z�\�{��+4Wd�Ǹ5�PM!�DUs��5f{��;� 'i��f�If� �����A=Q�#tۅ�<&̊�W��#q6�k�*���(
�)��!�xE�p���捭��{<C��c�Be��CLlIv�{��c��vW��S,�f��|V)TUY��q�8T� @M	�?�ͼv&��4�>��{pHp�684��6�?�6�*V���# ���O&Ӫg&��K���c��=�L!��7�7Z�L�:��9��^�4#�w/�2��vB��7E�c���3�s�C�Ɛ�u?��/ñSϖS5Ñ��q'a�QH�
;0d�u�'T�1#v��/	,�ϯ{�@��J���O�TZ5b-n�=�S�x��pt/��Լ�@(���m�A'��Ҁ#�>I�F-9�#~4f����j�=��]f-F`������mk���}7�E�!���"jADk��9@^W�A���t�D��I��J�֕�"�G�yk��iq��f�� �8�68�qω��@X�SV(�Ω:J���Զ����s��YO������g��uݴ���'�����d0��1S8��T�t1\�b����?6��?����x� k�Ȗkn*~����֙}a�n �ٗ�Ç��,6�j "q6�gΐ@髵Ư4;f���؊�Yej�$���I�=���ҹ2Ydn<��m�n[���\ w��4��B
"
�T�s��,���˴#4�d��e��Ʈ׏�S�����
��<Qw�@�B���C�� ij�-i���}���
2��A��5�,_%D�+l���;��x]	����r��!H1ħ��+��+�(+�N�X�w`�ș!J�t�8������y�c�F�u@����aۢ�c�(g����Щ.��:�`�����Ǵ�*T�P�-m6�
>P�$�`U[:�O'�ǈ�5�U�%6'�li��;`Ͷ���IS1n��9$m^\�0L�b�/'L�����bu���y[��B\��v��D��>@�k	�a���v���C�t�����4pf��o�mPȩg�m,�cbDA:��n�F�j+��5\cƽ�����F��#u�	���=\9,O3��b�u�R����v�Sh�c��[`i��%W��Qw�����mU�5��F�9�4Z�Ҭ1e��e�����!^�8y|��"�sͤz���	8�w��?�3rĺ>���`�N@XA�+<�c���lRMk��z���-�dWKU�H���FB�m�;�Q�.l�^q��ƛ�Z�/]<�4ah��{�n�xtP��g�x+v�Վ*v�Y(�pǱ�$��(ZLY,�Znrn���t����<9S"��x�Z�bh!��?nO���㕀
T��~);��(����^H!ٚW}�ٶ�S�p���ǈ8�Ն�m٣*=U��i��H-tS2H������-�w�Нn��O���1C���i�`"��� R!H�
��D�`na��d{�#}�mAn�̫51�r�����o�c�pЫaC&g�]��)��"|�覑�~�t��4���ĩ��<�.=��>����#6&��_	��&��%՝"a�wƀ̴S�͐e����$��c�j�n��H��Tj���L���73[Ɛ�P0��lc��{���E~�+�A�a��u��qWv��WH���bN�Uˮ�[��4�ܿ�H�QAQ���}�ʊ��%���H�~A!�-'ɻ�:(V���4DrP�x�ia�(��ʳ����	���cVc����g�[Z�cE�\�v���9H����M>=i/T�I�nx�/􂬑�^��Z��1'!����כ��Q�^�5LH�Yx�~��)�I�%i���fR��2��/&��c3��X�&E:)N�bc�@نD��β�����,Z-.|�Ȁ���Ż����т�mMh��q�kˬ:�}�>2�B�jY��yhn��V��� �Kw'�O
�߫ú�P@ߊ�"$���4��p%ճ]�m#k9�jRk��@��T,��"P�{7`(��-CE��lq�݉`,��c*39�ת�=0�+���p�T�����v��@��\�;.r{�����;�
s�z���1�Ϻ�2�v�
w+�����֬�X�!+�fUE��:O�5�hJ'߬�/Ȉ�"R����Y�:��9�PM�a�j�G�_���,.�M�[�6��?c���?*g��$(�����OA%�����yǛlg�� �t�3d�#n���� �h���*1��^���'����m���q̦:z5O&ݎ	|�骒֭��ﴉ�!*�U���S5�ė,o��v�Qe}�����-2IV��/:=soT���:w?��.���ʋ���@��_Z)Lo��]UB-��9|X�5��za�n��F�W��