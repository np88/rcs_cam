XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��_�}Z��BH`;H��`:
٨��m��md��	��v��|Br(PzJ�"���A�:�YpZCB��k\�ף�ܮ�+v�k&}C�*�f2TIj�_��҆e|l�g'q�<_
��$�gf�|��k�y�i�s[u�pLS�s�#�;��9q��}�O��� �x�(���k
r���x���[&�u�I��`L�M�z����"o���w�浑H�;�s�F���X�,MK7��(���i%E�M�H��a�q1p����E4�)ĭk���^;��� R����IX$��J�xS�싰��Qxn3'�F���l� Ƥ�
���$=��i]z-�v*L�=.IT64<ߩ�{Ns]˷��L����"�@��ebg���S'�D\����'�a_Ji�&��yx��z[���z��̎�^Q��Q�yt7�	�oB���V�b�$�ui�}\���������({hL��n��A!ѭT"����J�u�$!�i�]��̫Շ��㢄��o�y���ǘ������H(ڎo)Z����x�Q>���q���9��F6��H}�o�H�ΩK��q�t?�lU��r���a�p�n�}��ަf��%v6�h��Qm4�ނ\M	��jc���C�����h}POD�!9�y�����O�F��Vp��6��+���r�n��X(g�X��=F��ݳ9=�AV &���H�R� m�1��U���2�!:�E�iC��n�N���~6J��ݣJN�s*V�+���r(��f� ��	XlxVHYEB    b8a6    1ac0���;���Iw^�!8S�xZc��T7z�T�bp{XB/���2`}�������%A3
�j�;��%	��3�����p+��{��~��$����"��˛o,��܁���nqq*�v�����
�k�+ȡ�jB 6A�#ap}�گ�Ҩ�,afK�\��(޲��dF���B�B۬�oy���Ћ�8WG���r�aH?�<�%t�.�!j��"cG�(�Y{L��&�Q���U�n�\c0kt��/�(��0�H꬙\�4� N�=Om;���=�JL���a282��[x��?U�$�w��>�x�q!�_�3,�2.��?����t��4�Z��A]� �)����~��L�~��y=!0�u�=�b��~�����~�
�M�<�/[�%�>���.�X�HH�2f�u3?��n�]C5n��Z���� �'��]D��4?:Su�I���G�1t��ٍ$ �~����24I���("r�Tٰ̯�#��,R�[��ӿ�����aXߒUr�*]��D��a�f��I+E�h�]�V,_x������Y[�t�ᶘ[� �1.�Wϻ�1����@~mxX�cW��#+���	��~9W�d�0�?�(qM��a �ʐ�w,K�ǽ�TC����XrF�Rzv������h����PYY�`iB�Xgm,^]�~IM� ��|Kr�h-��� �'?	�^��������E>YJ�\�|���6tM:^vu�{ȮAg�������v�Y�st%�4�`��+�C+���uע���%�B	�ґIT%�&ǉ���ʴ��6T�[G"\k�#��ԣuC�H>8��C��j�h59��9�=$^���bRhZ�he�+�/���#'��-�y&��l�u���,�#��Dw�zM8��ß�4����z�@_,�����Yt��3:��׳T<���a,d���O��dl�-�7�u�L'5ݝ���=��d�\���w3k��,R<��)��V�{�8�z�2K��7�Cp|�"��������z�����xL���ةw�s���[.�ג����G�HO�R��}�D�(~v>�c�I�.ޥ�x6bf���-��m۶����D��y�� ϛ���u�Ν����A��m�b����)�&k	i$[FE��-��5�"`�pM�0y���M�$T���^��SZ�B�GCIK��2�N;�} ����Vg��M�a�¤sH�/U�S|W���K��mx�z�f\�͓ ;�����������'��� n����GM�W��N�9�&��}#E��V��d��U;'v��A;˸�V~D(�֋V���cRꉩ��F>c��jd�+�\�>:���qXǺq�33�Ö.��<Ѷ��ie��=�٨
����Tq9�G����g�|�W\ �v�WC�NP�����̙Y�H;�[�f�}͙�-���O��-7B3猿�T�5Ą�1T�f2gr7�}���ĝ̶�����NlB��ș��R��7��r�v�@�q8�~��1Ϗ�q��l��#g�JЁ����oE�ɀ��A�IJ�A;�e��E(h�:/��se��
"6����ec �,mD�i�T�Ffc��y�7�K�"��Ȍ��4�q�.?���A���j6�H.�>�p�U��M��5�Zf5T+�<x��l�g��#�vf�bjs偱�#�qr�3]]�+���.�~�ܾ��~H�n��u�W�764� �Gh��
+[�I�B:�U��-�,�}Ȣcd�0j��0�E?��]��������$�2\��P.՜��	`��3���V�>�z�FP����InI����S٘ˑ=���n��S��?8���T�!w�c8g�8��PPd��;\%=���H[���*�ZN�u�l�7ǟ��9Y��|�+k���ǌy<�X1h����'2��"��a�����{�,��%&�[5g���6��"��3܀�X9�(xGb�#�fjd#�j��5�E��(t`T!;�d_ڒ-+4�������D_͚���ng���;��_;M�)@s�v����cε\��A��4�~��^�"E���m�B�ߚ�G1�LA��X�c=I���DV
g�h)��-,Z�ګ�MT���a��<�í��ΐ�S����iځg��B"oX���V_ļ���z�K �h���1�䎘� ���3��}������Zѩ�3�1gnRJ_�c���q�K�����90�����x�����@o@&5yWMd�N�ݺgf��,�
g�Qqu�Y6��9b�"��e��k��)ҽ�'1r|*0�ZzBb1X���$H��Y��r�JPͣ�\��z�H�7%s o��V��S���� ��H��ȥq�ʬ@ue'�d��-94�9Gv�@Y��R��P�#�&�17#B����Al����`Jxܾ�b�:sQ����K�'Sޫ.�X��_��^�PmgZ<ټ��DvdZ�J􈵞p�]���ZY�oV���S>������[CV���Ɂ[`�C���7zb����6&$l�?�Ӽ�;���퐎 ��"UN���^%?�J�\��?/�O&z�E�6�?!U�
e֝������˕S}B�(
OBfa2��t�h���ة��^���b�J0����ߒ�0�>��Xj�-a���X���b�V���F�-� �b�%i��N\�fU�o�@S�ٔ:Eř!��%���X�#b�d��8���9aw�;�j��r�=�����ʻ|��ѵ� ���K���a/�N��p�d��z#-�wS�e��.�5��E)4y�����2���v�F�8'����K&R��4ؙ���*� .�Ȑ#zo������~��F�q ��߰`%�n�s����e��9|�m>��ºE�1�nD���ϲ��n
D�+����P�q�H�]��|���=�:�L����j2�W�;J犨u� ��n⾨	^�%Ρ�%Vk��-L�b�L֜}���˪d�r�6r�(�X9�[���j���$:�z)N���8��i�e���f����n#�k�.D�F��1j��/��]�䩚@�Cv=�gM����Ta>�֢CX�ɍ�@�HP5�pTZ*
[��
��ނ����/�V���)n�!�?ڈ��5�h��cE@��b�=��8$@�2�S��M��x&���4YH|1.���ڣo��OI�Ȗ(��� � WO�������C>���VC8+��1#��(w��2$C{�}}V�t�\hG�U���ے&X���.Z y>R��{�",-l*�À�h����Ө��ch$����xA�}D��r8OPCd����(�n�]V)�v�C �"��۰Vc"xΚ�S�����ZL�Z�{�|�q�5�R[���� ���G"�@�fnc�ۦ���'�G�j8�jČ��MS��_^�1^v�%C��p$0r���p�˯�����|x��G�2�	@R����Y��!�"[W�F-SJ�e}7� ϣ$�aH���V����^gP� �Z�����i?�e��V�t�[��8���J�Ő�kg4_d�f��cE�&��������qO�yn�8��
��֫7K� Ĝ����7Vx9�q|LJ������W;�� e>gGN?�;�ǎ���VfA0i�M���`d�s�ؗzU҃�
g�5�~H��Ԡ���p�P�V=����w�)�$Fy[ZQ���⎕�M|s��>.|�_�;�/����SeH��#g�)}�M�������42���:�����5F29��&[B>e;R��Y��Gj��K�$!��c��K	[鹣���q�;m"��u��w�Qa��^v��3C?p��ZJ��J��]>�EJ�ۅl9��<Ce�RK�㛪�KQE
2�,�\2~��nfb;D��l�Plܩ��$�J���@�뜯�&��BJ������&����v2��lA�8m���r���1����q䷗�	�<d�����1A0?�
�K-`Dz'���߯�ǃ-��'q�~�q���?���!���*�)��Օ[��b�"2��q���_n�#n��sw��r�=��z$��H�!P�s<�>��94Pgπg�Z�l��GS ����fϮJ�G��Bo� �**��=��@T�DW��,v��J� Ļ��q�7Woʕ��O�;r=)+.yc�Q�&j�o��}��L���G����3q-H�8 ������AF��?�|"�ty�S��lÀіݤ	�]��c7�r#Z�,���s�a�Ś�s��㎇b6�,g����)"�v�QgC�w�>Qf�孢;�pw4W�2C���,A#!E����7��Y���Ë鲰�����y��#�w�g<�Btk�'ũ	i����\&�[o'��3�5���Ƥ���b���O���l��͌��ur#���q�&�?_ٜ$ç�,|�#;M�@�5��A_�h���k������p X����B����+�e�')4&�]�;W3�l�q��mmS�"	�Hz���D�c7BK������5�!��k��r�ș6�-9r�h` QD.��������z��?�q�'V���{�懪�8�[&&EV� $Q/�d=�����	��Ғ�r9�ͳ:�p�	��R��=���I:��H�S�d��NP[�IO6n�#o�R��N��l���O���,-�#dC(P�[0�gQ[���؂�YPє(O����?���ϰbZـ���O	��ۧ��47Rj���vi���孭w��DG
 �H-��ٕ����!k4̛�;RU�+���|�6�T|b�ZR2�z��<
 ��?~�9직�LD�)�(K�%�Ɩ��i�k�l��i/`��=缄�J�k��`uiR.E�Һ�H�nx�Mf���MiQ��4�4�u�wniK��fl����Ete����]��/_�]��7K��D㐽U��d"�k+�m�7:&Ý�Y �t	�ْ�L*�T����O?"����\Ƿ�m�'j,AB�N[4�|F�q�p]4�aSc}җ� @����m���C����)j���GMTT��_����I]�D��j*���瞡z�����WG;��Ge�@<i�L9��UR�Gx[����幓#�����7�&�eK~�/H l�����`����T�7Q�RY�R{J��Y�o�m�,��<6���l+��G3�Ąʽ���R�ϕZ���>>�?�\C6�;���3=\~��-h,�i1=?9P+�����4��*T��4O�Y���,d��Z�T!�h9��������4|�:D(O��Ł_[Y1%�N�3d�F2>@D�C���rz��X;_$�iXFW� ���Z����{~g�^գ��q@
�_�u�CF	�����$
��!YM��=c��		�G�n]۶��6&o�����3l��I�٦�L�VV1���b)n�}�%��D��*�g̜Au>�\B*s���Q<�����������7iG�C������G��\:��t�삡}P��������*�mU��S��-}
����@3;F�B�a%����d�H�@)���߰�ސě�8i�a� OZZW4tSK�.�z���@�͹�p����<5�?Yɭ���֦c�E� r���|��I�,Nk@'��I7U)Ֆ�KOm��1�Zܷ�[VI5�֛u� g��#yT���@\����s����'|���$����>%J�#�N�"���YU�A����=�)�_L�mN��%�x~�Fe !F�������0��0#���*�޿Z�;mAf$�����ݩ�����#W�+��c[r�S9v��.�L�$���L�Y0/._�ʝP�G��Be�vH��g����<�*����^�1D=�$w����CA��۹�b�����ж䈶foR�-����Y
��+�Ȁ��wb%����\�@�w��T����8��Z-J���Z�fL�&�%��/��d7 ������O�O��h�dBTU��l#�9�%����� �i��҃}�.{���K�8�9���\oџ%�] .��c�<и
�����L�|��]��Տ�:���-�J���Vc$����|�نllq���u>Đ���Ok{Gf�?Eu'!z�U����kv��n԰I�Nt��!���G]sQs��Nf�k���utJa0���@�����Aɾ?"���i�]���8?��K=��JRx����f���\����~1z>V��-�j��Xv�f���fhRV} +R83a@V��1���U/�_L	i 䮴4�}X"��� ���	\CԷ�N��0֘PC���~>����Su�3��u@0��`����}�  ^��0��������8��Uh�fl�F%Ȃ�� =�j]
.!
�+,u�h�x9i(=��G@��<s��O��$bs��?D����Z3���nH�a	�IWY��-'$��I�_���~yz�ɖ|��ER��j���Lk���-����uh�1�0U�w�x:
�B޾ҭ�-O��3�����>��No�����X�Oi%F�5�*/��[c�����S�R��2�GH0�~�ғW�O\#`�n������?F�J�[��	q��M�t�ɢ�vV���ޙ[�Ԙ`�"fК�k�Z[�n$5=�&+�%�א���o4`o���'2|��u2�jM���3
ĠM!ʤ[�,��nWh$�Fuu�[�;ǢV��y�~ʐ���Gm� ���H��ίY��a?��n�w����[�m�����WI��������J��1�o��