XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���!$�`e��܉�k|���]Y������EW�[y�\����J-e`���>Z�k֝�P�5��X���D.s�]�q�z��������U�L�r�À z�� ��9�{��N.ao��^GuHvdr<-9�>g�Tn��f�ӑ������^鏙���YG�1�d��Vt�nm�������Xi��s�8��&8�SBWT(��/ǻ:��^lIP^���9}=rkLg�q� k�J�w���0кK�<���Ҟ�����-4��b�B�2�B�-8�(�<��T��V^���Q^�b`%S�7}y|5ջ�0R�z{ �'R�j��A�ݰ)$����Oq�4�>(��n��Q�Z�9I_,K3���)N�m��[R1Hy��ʀR���@�Ѭ�F�����A�l*�#6�dTsA�r��kh���L�T�����iN`fe��y?\�s�z��V�<�aj�]��+�L����ЛM4?S�.i�H0/Nx�xM��4�f����B��ˢ�+���M�	�e�*�Q�8�+�D���x��B�n�U�îR�9�#*�4��MN0y�xc���/*SIX7�P]��m`��!? ��F�����.�Jo��z{:z�AY��lG$�05x���TK�6�A�f��5
E[�BP������s҇�`�u��|ͨ��v��и��C�����1ۛ�4�`�b����;�EM��6����TO;�� E���d�oo$�bG�b�t-�t���I�$�U�VQ��������:d�r|XlxVHYEB    33cc     da0�w�̮d97w���5c�L ���q9uH��S�^�\�A:lV��!te����l�O��$e�_��w;x!z��q�o����+�ݟ����}�8aC)7\i0f���,��35��	j���d����<��Jٹ!&��]:���I��۹St:��M'ѓF􊢔�ܤK��x���ҩ�����Z.�ѓl�ś,���rpm,��\�@� ��ϥ=���$䝛�g���t�Su�vSTG����gH�Y�w�� PP���Ȧ�ۀш9�φ�Q�F�쩩��$ R�w�I�&��P���!9�
�ĩ�)I}z	&O�JŽĿ�������I2�n�'\0�]��B�wR3SW��8�D�~v.��-hxuqu�q[ysM���D�ς(4�ˈYs<���1r�ɘ�̂�N�]�w�ay��q2�=:t�Jv1�緜�V>����\��Ĝ$*?)�����'����KL���Dq`�[�b1�gx[� ����.%mMX|��b����A�c�����7F`Y���9Bi�= ��e=Bk��D�Q݂Ǳ��:^Hv�`�u�l��W�?jr�c8<��� ���|��bB�����b���F2���T�����@��=E���=eF�O�4�阚%�n@�Sc����~�+���f��l�S �B���ƾ^ܣ��+���2��sn�?aԂ�_l�6���YI$�L���(��1jp���'�/1*��������YȉK���i��uF�;�i%��d��7�;�H��PÌ��sY�f��M�0 <}�fL;, -C&���bS=�kGh�u��%���p ��q�$¿�On�S�b9꧕q��c�_��oh�᷒�����n����9�5b�����n�|��f�P%T$\���������0��{]�z���eu�fjX^׳��}�k�T(+ѯh�LL��VΨ=4����˓mLU8�Sfx1a�RT��(��;�������� �h��X��<@t�H�y%t@�Gʳ���㕺�_!�'�a)3;U�� ��&�{�����f)i\��|����S���z$����]N�����m���*H����@1t�4ɘǟQ��jI~�1�7~"��</��8/m���h��5:#"qskG���>X@�}�6�Q���}�����9?��e�.��f��R#D/�^��2��1��;�S�������]ky���A5ce[�ʙht�Bc���Ъ��Ef�<eq;��
7�0_�R9 �[S���-���v���0.
ah�
��+� l=Y�L,'K#8��Q��_qx�Z�
.�5���?Q�}_�!��[���3�P�)�n/<~#D��K����~V�$��~)XP�1���x=)�e�h��e.���\f�s<�@}[Z� &r5��EO����D
xz�eR��q���o�qt�+��VARt�$��g�maE�N
���Z띩r�b�� ?J��_���ϧ=��b���6t���_:�,O3s��ԑ����2�fgb&F5����׉^�b@�[�2\��EV��)xxx��!.��
h�r��b����ͤXM���q��а�,!�$Y="M\�HM����z@&����R��yf�+�7k��;sD�cs��%���5�q;��.���?�.ֽ���v�V��3�{+��~&�o�	o4�2#:pH�<�a��	�x7��ߌ��-n�NƩ���[�\��U@��%��ֳ���.�5���g'��x̰mIiU�z�X^�W�g��['�����i�8�8���gfT�*�+�	k.��y�CnRl�m[��Z�#�3��lu
����n�����LΦ�6���{�[G�[����W�x!���y�,�9P)z<h���
��L�Y��նT��/`�V��i��b�$E@��7�64���ܞ 0�1���/��F�4'D�J'ֵ�4��Fm���Eq�V��#\�Å 
� ^�O$�ys+@����ͺ-��(4�X��KX�|R�A��W��KN�V�:�ihvղ��	�X+3v]��l�)�r萔�
�xk�w����U�{�	_&�0d;!�D{�e�7�-�ՅX��@"<5�2:�e�=�����e�,0S����0y���6!�I/��d^�9��nt	�G��0�x�ߤ$�Y�*����/��h|g�6D�tY!M�@�!�E���!*���3�i���T�� %�<����%�m� ��L`zOG82��Z�������(H7'�+a����4�X���"ׅ1��q%���7e�n���dL�l/��w�Yg:r��ŭ�e��P5VP�P`9d����h3���ݷ��L2�S #6����e˽{	P�i�3�yi[��>��2���O�r���l�M�	gwU_���=��jEx��j��\������#	w��ڸ	�\q&m5��UIJ��:�]>��$��0�k_��d{�̣�y�7��_��H��6��`�4���?�1�m��#�K�����3��7b��Q�\`��#���!̦���N�ϥ"Ϋ���1z�v�%tT�'XV�i V`�"8��UT���ndbf3''���+P1Co�0G�N�2�Ҷ�\��a%�َ�2޼��4~I�kP�h3�wa\y�'�ɺ ��x�t�Zw�KT�D�/,�q�)9ӱ��n;�3��
u�z��^�@o�^�Gqx|����6���i������v{V"w	����6���1c1�njA<ه!�E����~� j/��X1Q�M4?��n���ޙ��;^8L���r0I-|l�.����� ����X���"�%H�랯h:R���+"wWd̬f
���칵9��|�<��3H�n�P��g)>%�ouK��F��PS�ҍ2sv����!�3�z�$t5��nɊ���T���)�b_g����]g�|p�	�z�6I�MT���O"	@�^J��1�v�X���N���H�n�
��2�f����n��g2��G�:�ȇX��h���<o~��Y~�/�/���rH��<.y�7��*�z�d���o�ϴ��r�e�������f\$Hͧr��(NR�6��6=�8�J7��>(�nt1�1�v�Kl��Ѿ��B�;��;D>5�[�*"�@�V�Z����eu��^,xON�)���>:��lh�j"a�nk4�=� �7~�ǩ[k fb���`�ʓ��|O�|R��w�@@b�>`�`�G�>�] ���*�_�y��1w2�R�V�
��e�&�i�̊�<���#9�2�����H�
I|܂N.�z}��b�c��%�h���&���6�1	��������8�߈�u:��-�
C/�B���:	�\0�������կt�s
��D+P�T-���T	2z�R�%�D[����a�]z3��{�pR����<m�CH�O��e�&RK�NF=eY�:�Y{��p���