XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���Y#���~+ʥ�_�,MQg�%݋�S��C����B|����2�Ч5��a��=��wnQA�u5��w�ׇm>����p�Uv��z;�����ҫG��M������G1ӏd�ȶ�Y�3��U���S����ac�c�֭=�x��˅�ɏT�`/I�B�DB9Sf��g�Bm���$�</�������S4�	�!2#2�*+?��c��#�M��S�����Z�onΆ-U��<�J���`&k#�W'W ��2^���Ƴ�w����!)�&�'���ǳ�Z%�hF�doEd�\���� �������P�!_3^�6������D����f���	y���(�ֽ5��p)�AJ��-�p�����#�Qj��I��%pE��
�5����b`��� r�aO�r���;f*�b��~���(U���)-OZ�R��}�	��+�k/ �a��socc��!��~��)?�(�W�G/5�$�|͑��w ��w�r,�0��=݈��F=�:�B���8�Iy��~q\Wp����}�;і�q�
`��������>�_X��0OJ�����喊�C����?��؟O��_J�M��K�ۜ+��dPwNΓ����Ss2xVɟOS���ͮ�f:��y��I���f��)�����-ʍ��F�����VDb�1nDmE�L3����Nh]���!�b�S���s��~n��v�������T����a��wG��F�#Xm��˵���n���0�XlxVHYEB    fa00    1790:5A8���%�.s�
�a���16XK2��¶v���{�@[��Sa��.���i�S�k�p~�)�>�TFb7�X*b���w�  ���R^�n�eaBK%�n���F�xʤ!��T	�|m�������uS�δ��akMpm=���N K�1�d'7<'�����>�ݴ�ߊ��^(`�W����Y6]���Oci���?-��}gQ ��)���x��f��&��E��e�E.�$���G�Ӧi��p���*��*�P��}-$�/K���{1dPq�L:mC��j
�
M"�t�?�8%? ��s�c�4�Е����Mx4̓�a|��?%�,�ۏ��7�B�)ӎF�ί�L!�<�!�h�^��27��b��_&�;^��]��>D���j���uZh��(���=}6��-I9�g������Ehn���[/_
���ߤ3�A}�����cW6�����mv��y�u��S�X>�o�\�����Gjc�[潈�y�-��^p(�a�J�_ �,����'U;@���G[�8���"|��Xxص��v��G��Զ��*�Qo|ޙ�GK�Y�����[Ƌ�=!�_&Z��acQ
���7ǃ`���Ģ�,��Ѻ��%�u;�3:�|10HA��+N~�KU��'\4g<ʕ�*���{��]�R+�ǃ���Aڣ�T&�);iC=7M"?�y�֎U�w�Kw|�Jø�8e ~��PSY���C�ˇ�|��L[j� ��Qʟ�"v���G���~a_��,&HF�1˹2����20ǼU[�F)�sNT!�j��T�}��d�E�`�X�rN��R��2�+���B�e�B3��d�v��|�$���s�m
W���:��
8�X
�թv~�k���۲��L��?�Z��J���CZ�A���[k���.)�ྣ��gytC-)J�X�Qr�o�g-·�Am'1�	EȪ>�>����H�e��~��/�6f$��	E�,z����D����lUT���L�2�ȧPigOG9�����7�NV��lIy�0e�n��8�2�n�T`k*��4��9
L8rn[�E�B����Q�NCb��Xߜ�t��!5������ӊ��}�H����'��z����z�^��gjb\C�X:���Z<
�65�n\wz�Y�M��(�t�k_,�F��g�K��� �/v��*�ߕ^��I�6�.*�H1�4Qq�׉�OɚX���2Aw��\N�ʰ�t`�% ����|p,���@ݗ�=�(O\�U�(Fײ$�ꅊZ�p�;��M�etvV�:�:��=~eʃ��r9���礛C4sl�p�P�7lv,o��R�.�:���,u���p�{+}j5���x<��o�;ke*�}����`�g3/悇��m�.��*�~�o���D�ݷ�d�I���z�љ����d�	�ǁ�!��P.����x
�^�i���{���B��^�����n�-�iKe�+���"�1gn(��/Z%~|�5c�>O���#m`q��&�=��SPT�\���E0L���J_iZ��N���]����I�R���'�z��� {��y�!<�7��b������l���l3�[5γ�n~�v~Z���,$R������_�%{[W\o��%�T��V8�]��Eܦ�5�)�X�-JK;6�70�q��V\m��-�"��
H������H�X#�^��7����X��ě-�OT:�P�_��\|ق�����3$k<#Cď9�l� �qhO��aB��r���-Q��rxS1^���2�c6>�k������G9�baE���/��g!Q�Rl�wu�����%��֚�d�����tO�~��|��VJ�J@S��i3Ǭ�ɫҚ��~Չ���@/~y�$`��=Fm�_hX�E���	y	��9Z�C����L���h���_�'�����^�pgܲ������S�V����4pcS�l�H&3��c	UA��y����\Po�u ?��VU�U�>�y�Fah�Da�q�H#�S�W���,k����v�>����ҧ,G�}��7���߅;�G�j^� �A��wx�ƞh(�T��Dh�h�T���jGJ `� �����+����#)I�k6����;ꮵ=��>�mm&B�]L��֭���j2b��
���]�P칉UF�[������dm�����1zn}j,��D�F��uh���~�1r�d��U���^��SL�)��d��X�+�#��m�;d�����Z�7���u	T��3���E�@���_�9�\����"2	C�E&6� �bǯ-�D}Gz���41Nx�e(j5Uw��|�/ԅ)��PА����܈�{�lm/.F�����0d��_-��H0��=tK�m�U/v��w#% -?I���'
4��ͪ"ʲ�Ds	�����.���!ɠm��̼�S���nX���B��lP��yN��O%e�=�U5��kr�#��'�|�I/;AAle�w��^̈�=�� w=�x;hj˳	ψ_%-@YWDܫ�O*�[F�G>�Uf��1m�J�>�p7n���vQ�o��ћ�,���hXsw �r��%��ͷ)�_6)��{d*:��b ���^�Xb��b��D$G��f�i+���q�}�Y"*c��n���KK�-�%9Zt����A-b��,�Q���eDr���+���������*�b��g���V���oj�F�{ӷ�ȴO9Z�����	����Y�R�@�<�QU���a	s���Ǘ���[wYFv�$ۜg�*>i�jҏm OmK5�c��6�d�����YZX��P�a�ÌMP�2պ�D_E@**�I�u�]K�lD��H*�7A���s/#�o5�w_I�(~�늵�=�#4���PD��/�o��j?�ǐ3gO�q6��~���V�^b3�K�Q�'r��5ȃZBdE{�<+N(����HO�f;�?M@��+=0�8m�6M��s�Ry���e�� �q%M�����a=^�΍���]��:sZFM��جܹ	4�m�U?(��5X�(��N�p �S�C�v����n��Lt`(�<�}���Ÿ1R�C��<�*#0q�S�O�B� Qt��;Rʋ`cL���إ�����(r7��k��톼�[rf���9�ș}cn,C�J�Pp����ٶ���Z��\w>O��XL%^r�8~ku�(�}��� ����58�p��w)|x{�/�PU9?\�R�/��n7��>]W���xg��0̨��f��@^NNX�Ȱ�̦�>A#�7n�>P�����ayeZ�7��C���_9����F��5%J[��N���[<-'mMÛ��1�t�ݏa^5#L*H{�~i��"��q�};/Ãdnze{ ��آ��\�ۙSw�w�Ɂ���FGq�&_qr&)T�;0�l@`�y�\%�d�G�w�d�z|�*�Ȍ��DC~2W�����n��ܰ�=����f��.[+����U�tT�!��&b?P��*��s�H}-=d�]���2���^᪷�a��>�FZHe�l���؏���B���:���?"5z�kܕ5c�?4��*��*�w]i[�	��Ky�>�M��},�,D�E;�f[��e�����N"�Al���W
������	�!��7"y���ܒ&�;
굼�������Seo$���Ƿ 넍y}����tr�P���: ۶	� z�Z*��.5�U.h��b���'YHm�+�uޢt�O^OvI�*o�0���PI�7�+���S�l�Ĺf�)�XS�D,H+�s!9pY�������;��wO���偳�O\����'4>���!�\N��A�i��zQ���E%O��^a��}LK��燃ϯ�9�ַߎ=����o� )�1�3nE�/Edt���ck�'�$Q��;���"⁠j�F����Ý8�QC8�T������4(�����i
�:_JB����x��Ԕ���S�;�j��Al��~�()ދ�<#c��*�g��2�����E�����,H�o��@Ue����A��t���T��gI�(*���L�����=(z)�˪���> ?�WԈ旓|<� �=C�%��"��黒�㍡J�P�a��ͤ�*�ѳ,Q����v�tB��Ћ�d�. �Vi[�>���P�����Uۼȱ�ю�]-s�ϧ�̟���аP�'O(��G���*`�ۥ$iu?�{���i�#��d0qr����y�o��p��o�᱄�w&d�A��a���Q��&qQ�����"����q_=q9}'��t�=H�=Ô]�+��X\��;ĝNP�f��C[�$G�@�62��2���ߟ>[e(iA3�`��<���V�f�PN��:���f��I��C�/X���/��)�&�/�K��bQ���Ge��k�$��sABw��)�[��nPV�Ҵ�}�,���g:���|K����H]�A�ӌ*#
�Wl�������fg�����`�3L��p�@��:8|��d��f~xdbZ����� 3��Ȁ�_H:Qq�49f�A��
5����nHy�G��vѶE��4��F�����iL�`�#P&�׎I���f{1�W]:񊤂�����Z�Vt/�bi���/��Fe�ma+��8�|��$����X�-�Z��^����K�kb<F���L�&For,��SQaC�"Y�g���U)J�9ߥQ>��\q� ��5{�;�l��O�����}����0n�2��5�4��2+���<�k��'!��?ӂO] �*?Ѻs�*�xp&�/���$%C����c������F\_�@<�Uq�qy�g5��
��o�No��J�o�$J���ׄ�w�Ў ��Y�pF�V�f����p����)��a��c�=Q�ŷ!��(�&��#d���=������!|v��7�Oِ��6���h$R&j�A�^	`�Ϟӊ��Vu�3�,UL�mG8�����,�'�Фz\��yv ��rG���G��yZ� �E�xAj����T:fn'c= �a��T�Sc�yx�I�Q���ǆ���f���ӊ7�\F�A6�i
*�_ХI��`Ѹ�����u�������g;g�Fek02�l��mد+"��,� �<EK�'�r�j"U��ڬlЩ�J�b�b�e"()�l�n�Âݓy��9��������'P�eG���,'9N���)��G���r��*� �*��O��a|��s̓(�Z��n��e�2T��S����?�i��.�o��A}�f�0��3��E�������y����R���DΖz�1�))����6c(�խ��?���8}�8!�6�!�2W+�����W�N�۴T��U)�cq��6�x�m����z�	BI$��� ��K��J�I�{bz�j�����'j�m�Pt]KPjB�ZS��*�� 3��	�EQ���A�1�ú϶��\Z�Ytv �9�{����xV��?d?���O��n�0m�g��#Q���ir��4$�v�V��A?�2M���Sf�N�q� ��@����e�������##,�Q�R��N���9��[��H��훊a�L��~?1��O����'���T��v�]j���uU�:�Kl*����<T��k�U q�Н��U��n��y��)8�)N���N����.,���cr�A
���]�X�<'��Nn[��c�zmI
B���I.s�A֬D�C�B)a����1H�FG*�L�n���B]<�S~|`}�������JN��Z�0}FJ�-!lE.���ʣ%F!�S0J�w��%�Xդ�i�a��3�k��o�g�5��~:Љz���5�>���t���3H�u�1Y����#����eԶ�0.q���B��F���$��_H��(�*X�<�
�N�[\����]7(�_�GXlxVHYEB    fa00     5d0�򷎃���Z.pq}���2�`�1UE���T��nlb��n5���$�썖L�?���TW�N�1$إ�:���b�� �Aێ����4�f�Nh�Z�b��y�~y��~r,{�<S��pò��A-����j
Eq�� ���;M��Ƒ?\���uMcG�#"�ʬD����KK�~`�94�̢����^���R��o�i���oV]������1�vܻ��l�rn�C���M�����ӣ��g+v�Ė�<5�Z�PQ��,m�$-}?��f���WK�j�*@�˫Z��z]+���\,�1J�sl���w��i�"����#P� X�~�Dk_e������?��£޼�����	\�?@��7nzQ���-_�a�lt�\/�$6j����T��`2��� �����*n��&y�G+b�87�QD��!&x*����"3�4���)�x7�G��^��I� g��
J��������Z��lY ��zI��S�b��@ſ���q�)8I^v��g>�+�7���k�'��1�4�λF�_`� !���M���^ݐ�y�a�� ��#��h�쟉F>͌�-��Gљ�X[s�뀋[���H�.`���AQ-�K]�>�8����G������.]Q25������*�)�ˀ'vܢ���(@�Ȅl�P�)��vc�î��@������x�a��}�0�|AQ��}�����h>&<cz���Ʊc�a�a�����|b�������>$�+������UO��0��B���9��.8h�B	.Ϭ��N�o�����6�����	~���
uK�yz!)? �@����_Bsq�^s}F%��u͔{�p��(\޽�ZR��%H�I�`VQ]��x{#ix����	$�W��YN�
py��(�*��=�ʶI�|��ص�Պ -@@�*��_�!��p�G�/#S�*x����W�
p��������Z��wx�e:1���p����v^׋�Y_fb(�p��Q�(Bh> �B"�y��8<x�Y�j>�c/)썫�I���-�/9r�?X�L!ؾF�Z�榝�y�A���2��`��_�y�;ӟNvHn�����l� �3z�& �}Xv�W1��nj�󯯄��|a9����3�cC�r��HĈD5��V�E�.�D�����Ğĳ]K�8���E/�8�ۏ���/jKb�r�^����Z
>ԕ����s��O����{�'C�{�
������A��3�^��9`�/��w�_�p8���l� ����H�,�>W�xgm���%�g�KéU�w,��(p�3�7��&����[?I
&�n�M�wR�j����z�v�^��0`����+�8�,ۣ�OJś��� �T9�_r1�V�5��^HΕ�ɸJWPT�|PjT�ɋ($Y H��Kⶢ	�e8�}���|G�y��%��=c�u�71��Y���[��x�@��gF�B/|��#%���IXlxVHYEB    fa00     640f�� �!S7�M�S�f����L�X�x�8&�-9jS����v������.J@�nϽХ��Q3$��G�ʺiz�䯆φ;�<�Ѿ��V�;��8��ԁ#�"E��U��jZp*/����d]���������b��c�q�X6L��b
l]��B��5jE���^^����Y5^e<��j�c|C�P&��A�+c�u� O轱�ͭ�e>���O��փ��M�Qc��M���4���g8μ?
=1�����oeãa;���n��q��&�֌����c[��k!h�oLS�ǁD��t����+�5���l�T���`�AK�9���T7���n�� �.fֆ�wQ*7�N�J�F	P�g�`�D͏g#�{Q�ZaɿZ���q3uJɏJ1cF��P�F��C�L)�p�����c>��o�]n��w}N��N��p�6�N��w�v܆� �@7��=O�7�'��[,a|$��A�HՁl����ֲ� ʄ$�z�x���Й;���A�#�Fx�=�hn�����]sNI�F������] a{2T�ߑ�5�fx���bD�<�i������x���0�����h �h	0�)z��a�e�H)����ՍVkE�q^��7��(G��i����I�[oY1�^��_��>f6�!�3�iG�|G�/���&�t�V�&������_.��J��q*��N�Ȯ��DqRxe��=�N�8�P���Ar�'�آPu�����Mn�g���HR����?�p�(�CmXj�*k�	���k��UI2�ѭ�57F��@g�s����nn�Ir
��M�!Q 1�8�L�7��*0����i���1ʈ���Rt1�]�Dn�l"Qmкl| y��|i"�nlX���pI�rƼ>����¹#��)����Y�7�/��:vj�r+�����ˠ������^2!�T`��^7��rՀW8p3G��Pe�OhkD�Eo����q66�.X�����u�+�$��Ch|d&�o��bp�v��^{��>�W��ux�T4��>�[Ӟ�У�c�Z5�ߒ�x�M����j��6���c�b�I��e�ܙL���떤oeo����t�����P]Beϸl��h/����q[n�M�-}��;����f;|�����Km�҆7M��@?0 r	?�t��9���]�`�<�֡ ��Re��p��}��X�x�Ov��5�l�oy;e�˓w���.�U{ّ��ڂA�bZ�rFfUv8�[�kM�_��nzn98��~�����	�yP�k��)����"'�.��	���`�����ޞ�	ڱ-/�񐶎$,��F��[�`U��#~�p�Z���l��z�ٲ���)v6�hÚ�����[��T|���N 2��j�:1y�h��c�R���`�2��#�hVx�� �zA�*�|��@ܺ�&ؑ��$��N�]�W�cp7�����6a��(�zFg�ɀ�7����z�b�C<�_�G�ķ�B�m�Ʃ��o��o����͒V�M����Z#)L�V=�E㙴-��s��M���Z����S�&�9�p�XlxVHYEB    fa00     5c0m��T\뙗�{{ߋ;�G7��?�D�����3h�+��CN]��0h�Àɟ}g>��צ�]c�Pr�:��e��D��"�k�"�K��_e���8g1���y�H�;��&������sC� k{�'�ot&&v��W˵�
�Z�sx�O��b!��u���h(( ��Ĭ5F��m�rj���P�
HTb�$δ5��@3�&�1�Zabu}���E�g�c70����aR�� �I�����:©��(�y	U)��!�p�[��z�:�͸�aD���w���S��	�e�{p����X�%��Zy���P��]z�iug�_�T73�5�r=����35ӣ����L~�>���u�oXٿ`A+����}��\G-���JA�YCP�o,�<���_>Y��(I���5�zE%��3�M�s��V���S(;��n��l�z��XE��L�/�F�Z���n��˱�`{���K�7�|� ���=���}���`T����i���IɌ �o|��h��v�&�����4�V������������7�8� b�@���9[_�J�� M/*�F���$F��V�f%��"��^L?�z����գ����ط��'��32z0��0��x������0�j*_�JG<�R�_j�7N�0�>*XEgt߱��{ �L@���,^zJ�BѮ�n�������A<Љ������6HV��#{Ȱ׈���s��WL�8^f��e~эg��1a��2|�4(8`H4ˈJ{�p!��1�L9yTB�vx¼���X<��G�qҏ�nK��N�Z[Y(9W��	�q"-��z�P���Ie���x�~�������25\����"�x�`�Tu�܎M��_%�q����'-�E!�+v��Ů�^�)]��¸���x?�-⍀�C$��cK=(b�_�Ë ����Z���g��������
n{}�͐��>(���S#��'YHo5x���q��+s��l7 "��&����Dh����ؖ�͝�^0���n57���j[�F%g��@�P;^������Y�����y_�(�����^�O�C㩈�O5Y�a���b�?,M洚LK��*�1͔�w;�6O��r�c(���E |�R=�3����`M�W��$	�:9~0�J-'>�F�}�Tv��Y����g��.0T�+}�Ź�7CpS�J��5Y��M#���يָTRN��r �,K�9�Mh�k�Z+�t�NR�k�6Zn#�y�����m��w� �ڞ;O�F��UȈ�L��t;�ݐ(#�<&@�3�%�1@)�u�h��T�8��sq�mhRW��]�	.��yg`�7���1�ʬU�V_���T��F�������&���Z���������h��L:	˓@</�}i��z���~�5�w����@���=U��GL=�X$9�R2�ᔇT~��l��b��� ��B�#�=K�Z_�XlxVHYEB    d347     a90F"��$��^h�PM�Gei�W{��9�[s-F�A��k�l���ԁ�7��ޖ�1b�~�ޣ����ȫ����\�fa;�rx3?򞙋�k!��ؼ:-��F��6���(��~�\��Gu��I�2"�ɇ��wxv�}���t�~��;�E�]zJxiU;��&"���.]��q6�gY&�8�v��NQ|������ax1��I&����n��@��x,]HCf�#V�۪�Gs4������gՂ�E��a<�gՁ�0��=���c�x��V��?���s�O��y[����x6�\����U�l�'1���'���X��s�&�7f�Ǟ���X!mP �y-����7�܋�!i���)����`4|cA��G4�Vv��"�l���3��:�5�(?�"C�r��o*5�e/R_�N�`�'��Z�j�,LOKW�w�l��DjK0���� ��c��,��h�kTc��}�&�ez��p�F]�#�~�~�)F�N���M��c��9�������M�X�1���Nm�.��� +���
��
��d	�1��$���kM��~T:h��CW- g��V���]u����
vCK��������mryI�	Wؘb���w�����qmP���ο��_A|�&]m����C/4o��"���,�A/o͓	r[�ar�z��'��q �9K�����@�`K
�6�b�q���H��l�]#_ъ�T�9�Rw�H���FX� B��fG�s��f5��}������:���Hkn"k	�z4�&WІ]V0��V�&��>�����u�drVU�^�=���<�eWxXN^�	�Q�G1��_/�F�;��|����ܷ�㯍�boxR��l�%]S�x��Z�a�1co�ok����D��i��X�3$�׼,e�+��T��pC�����$n�y=�z��8)��\����idP\�Y�L�G:�,:8@͋w<���;_w��fN�71Z�eT�U
l0J	�6�xy7���D}��3p$�\�|!�'���6�J�J{�5��t�5���Rۅ���"���]�7m}R���I�K{�J�b/��WM��6�ḅmS)?�y���]������ٕ��#m�:�x�bJ\�9�eF��U���R�u�8������,�d���L�O��!k[)��ޢ@S����h�@t s����D�J&��%�i{7�R���6�u�T�'��������HFB��G�դPGLy��^3�9�aD��k$e>�����e�+�$�v8�*�ٰR_]�b62��}���v�Cy��N�C_���%�K��_�D���~gh<y�<Θ�e���f��Gx���a�+�ͣ��T�d�*�^�������Z��L�G� � ����j���k>H����:k �$�`ݛ�&axO0����	Ⱥ��u�H=f4L��@�Ɍ�&���]}�Y`��q�W��Qw<�2I���Ru�Nh�Ai,�r����μ����ڠ�Y��URbh(\�} *ey�� ���&uӤ�S�֊�RZ&����`x�}�7r���`�d�H�GU\�7�}FRdk�m�P��_)�!�-P���C��;��i	��F�V�"��|-ai��pҀ��՛܀F��o�xcX\0�Y������\v������<&~$#��F�s�E+�W���r�tf��B����S�d���Қ�
/�:�<"*�H_Iښ����G�K�f_��4�J�{�P��Z��s��CU�I�r[|Z�Bu�Y��G�V�r����$���r-�y;�{�-�Z�FY)��4���E�?ZG����.V�b>xsk"a;d\~���!_�b��"\���R��,�K�7v�Z��D=@_Zз�	wi�{~�U>tZ{dj��0�?A c.g߮�0^�A����Ҿ�Z�U�Ͷ��5�Io9tr-�u�\�G�J��sK7xE+"��������1��3s?��kDn��{�+�r��GLq�	.YAbx�uO\�LLڛ9Xh��Z�� �A�!N�O�K0sg�&E�JX�u����}g�])��0�Qd#�{>� �}�ޜ���Rv}�GȇwG�mTUJ�	��bA��4N>�&_0�[��Ȕ�kxe��b^�=Mx*�x�+�	��Mg�R�K$碯ַ�wfQim�U&	�s8>12��z�����27D��T�,t��;Ф��$� �Z�l�D�7)���U�d{gͺ�S�����>��o�u|`p�*��bD��٬5�P��s���zj^Ө���F�z�"=�2f�X#�힋W���ly	+E"��3fՖ�^B%�Zlί>Y
����L`�e���@�4Z�.D��-���#����S�o�YFC:nA�kV:9�~�Mև��H�ˊ:��n�r��I���Z�����y����V������9�5�1�NUL�9��:d~���3@���i�cϱ�K:NRa4k�O�K���M���F��Z+�,����6/1��Rh�e�=K븑��E������vB��(���I.�A櫻�7�n�&���* o����B��$�蟢K��©w׹˥���I���n��G�>W��h��EV}�q��|ʤ��ӳ�_�D��g����/@�y���|p�N�Ș�f��|�_ę
M�1��'���䬀�z?