----------------------------------------------------------------------------------
-- Company: TUM - RCS
-- Engineer: Nadja Peters
-- 
-- Create Date:    17:21:59 07/31/2012 
-- Design Name: 
-- Module Name:    fifo_tl - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity fifo_tl is

end fifo_tl;

architecture Behavioral of fifo_tl is

begin


end Behavioral;

