XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���!9e+���'�W�2N�߇�n���x�A˃΢TG>]��~~�W�!oEQ��5�{�ޡ��q&Wo��]p�}Ah�ׅͫ�n�+�cd�Un��q�^��I�x�[h$�v�%DS7���� Z}N,Y+���X�:�e�89�I����Z�m���!e�n�]ē�MP�x���ϖ�Vi�#l�C(��}�,��c"�Y �!bq�ò�cIq�Vn����/H��+I<+$�j5�;�򭀜x�0�ƇX��f3�8�]87���%T�8�p���J
y�{�"ۤ�Xd�mQͿ�'[Mq��&7Y�s6nӒ���>��k�'�Jn~K�B�.J[��\�	��Z�<n�l�Uy��e�T&�sN A_o`9�`? ���/�d�KtY
�q]�LGTF �3U<����NnB%�<x�=��G��x�`�:�ӭE,��6.�d�+�q$��Ħ�8߷��y�(�F�7w����CVs�޽��k���n��4p�U��Y,pZ�����]m�0��|A��[��N_<<��d᧤����*���8{v=�
�품z�K��z��b���/%' ���I�;��c�H��yt�# �v돯�3���F��y̟��a"2]{)�:כ���a|u���nNM^��qU�t��V%�7�1$0{R�9�m�HH]�1��E=�@�)�v�x�������M�"<�!��
�ҘJ���?�ۤ�v��~�~��)~�� ��NS����ft)���$r�+��*|�T(��k����@M��(�XlxVHYEB    37dc     af0���+�F8������TA��X�e��9c����Pܹ�9B>�f�uK��x���,Lx�2���C��Yc�b��/������~� :�����;)ߑ��P���Ħ����4�H�ˀ;S���R�5�`�[���{>ɴUb��G��64�4�d�|�Ӭ��I���CL(��^��w1oC꣥���S��o?���f�E��0�V�'D�W�"L"A��A��z��B({U��u�Ϗ��jƩ���p�V��z�2؛G�0�^����];�;×��8�+ӧ �������qn�4ls������^��e������Ŀ�btf)��;�	&'��� U;�C�|��t)�L��b=+���]=���BD�}k��1d��#�<ަ`�5�3�V�-�����g��6Z��Oe��!Fxd̮�P�q�8���a���
���A@Tnk "�6c��e"�lE�sRm_�V�4�5K�@���F��kTk<$����!uR)gj�#]&�ɲ:���h�MA�h�
�
	n��I������d:a4y"(�&���\j��r�)r�gtJ0����:����~0�9~s�X�{�� ��l��9;9a����Sƽ��J5EF���7@YSؼ�]\�F�E$C��8�k
Y�U�$��5�1���XU���~�\8·t]M$]'����� ����٩J+8���O����%z�e�ﱗ��VCfu������W(6��m
�~��p�F-���]�N�]Xq�1�>:�6��Q׃ϴ$bb�Y6D�'S��"�c�S���$A�������>�_Y)?�	�}��x\��kD����
Hl!G��9�.����k����u�Wa݋��y��ұ��B4VY�����͖z�:�fC��<�!��L�y���&��������+��e��eR�F�Ț=(^���MYC��wE`��=�6�S��-o�������61]�W�*�@��1����|�C�� e�E����$���Zs�:t�����Lۚ^F!ߝs�|�%Zo��(�!xA01�N$v:ws��|����j=,�F�;QV[�@��� �wk�h#�2u*���H�ϣ�U��jj+���X�F�Dk��֔h>��7(X����<�k/����r�dh�b��{Ə���'W�$�d�#�)U�d�:i|i������Z��6����'Bs�d,��v�$"�e���=�;��ޑ�,�����"�,E6-[���i^Kc2���M�ɸ������yb!J������W+�y��c���O��4D`��"T9��G�C��n��͒ԑl��o�n�4�na)�'��u-VIy���Ie�4ނ�Ik��ma�m��П꧲&FXgPK��Su��'��e�A�ęNX^NoW"��D�A^��,���IuQ�"*�0�l�k������5m�ą%ó/�+�Y���4H�5�,�jS>����l�@��d��a&��Ӻ���E�)��(��J�
��L4���O�X_-�n���0� ��D-���@���t�ʡ)ϳf���\h����Z�9���,�5�v�BLJ��~�^���:&���e��e��f᪺۸	e��Wt79|*�Ll����:��K���t�&����EYltё�!ӌ���m���7+��>�JG��-���{�xy�A�A;	�����xmg(�erz��3���!�:�!H��Txi�D{u��� r��h����b^��#sv���i�rD�|��m���Z��~RY�?��h&�8�fK=�e��zZ��,?\{�u�������?���4���Gl�2�x&v�q�m��ڧu�n�{�����Av�Xβ���r�
yĶP������Pjwd��4�	��[x�������'B�R�}��-"��l-TY|�5�]���Uנ����0$8��z��N��
|�F^C�*,��T���VK�~_$��B�:����-踶P����r&�w�mr����G�|�GCC��N���b��`���@u^��̏�p����*��+l|��c���j�TV����Cɛ����_AP�C/9��B�P용�҇��D<fD��x27��������2���Y0�0�Z����Tya"+0�Pvd��Ž���N��sZq���$UR��y�>�?�o�g�����̍O��6{�����]_����hްakpr��AAe��>��'Apូ�O�6ۓr�w�y��W:Zc gR@����"%�F�ơe����ĤM��^��Q",�H�T����%{lF�R�jQZ�*C'�p���x!ˠ�I�>W~t���
7���-H��0�8m�m������:�=4�{?���R���̂QN�VC!,�0W�?���f��!µ`(�"�.~!�w��z���m>�~| �b�E�4��X ��9����l��Ķ���Zf>�� }��.z+!﴿�}�Ž������������Q�pSb'��p�S]DW�t��؟*�-j�Or�I�5�e�7׵M���|�}A���h��=P��p�φ6��L�<@�C�黳R�p=ȫN<)cf���xM������X3���K� .f�C^B�~rU���4�~ل��������@ouT$�Cln�X��\�)׹��O��M^���M1������Sd�_��g�R~dY�q�����3�u�g�C�دmU�L��YU=~qa�pM��z��T���Eʘ`�q��f�z>����[+��rqD���mor#���