XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��kp�x��p�}o�G�Pg�:�):�XHu�D��p����O&;o����5[�c����L�*sV. ѵμ��?��8�ng}��#V�M�#	�%\��}�is���������,�l6 �@���7~iC��D��ֲ�|��j�z�o���}_�r���fr*'P�s�,Oє��r;Is�+鶜�m�'�pX�Q�_�[�W�ߨ���lg��h�*������7x�R����kd���H+���C�)y�V{Q�G����������c�*r��)�Ʉ-<�[�:��Z�T@J4&����[��3)����.�/��[Z�'?�-�����f�g �W=җ:<�h�5.��	�,�u�y�me������Xμq{U���U���:^��+�veꗺ-Ls ҂%��9�`#��-� �*��$�Y��K_Xy]��:a2�Ŷ��K�vQ�4�AĶB�����."�0�l�^���bF�0����e�sc�Ah���q�`[V]�> :q�!��>��*SH�x�2$A�qA@��T�	�Ֆ�L�r)�>U��Bp��q�"���yUl]}S�R�2�q��(+j6�K�����H� >H�9�M�aJ
	>4�8�yp ��a2V��� ���,�,>�+3�=� ��j�
��j���(<��B��<!�l�
-���j�Z�. D������2^�L�W��%˰ǻ�Ac����,1��߭��K�����U%����q]�5{����ing^�)E��r����������}&����XlxVHYEB    9efe    1be0\g�֛#�0�� ���J&~�yOC9]�o42��"#��1����3G��wA��6V�ū{�����g�t<��?Iy�E��S��+���2��u%��&�n%���t߆.�R�P��Y�ި=s�|�k��N��vm�խ ����#� Z���������^��t*�f`�<��b�u��߽Y9ğ㚪�r���.�f���K��V�^�̑��q�̑��:�%o#�DuY\Ha�$Ǐ��kGG����`���IhL��B�ς$���������i��/�;��- �-˜�#V�Dnd�.l ���G �r�k�S%rE�W�d����.���+�i͛�Ĵ�fЭ;iuL�b^
a���mu���D��v˧�_1ٝ² u�� ��Z&s[U��n(���[H�@ߩ��c���,���c�L���͹P��ULN�6���D�pi��S{���¢�zz?��9��4*SGR
]�Ӥ�h�2�3�D��T����]w�"��E�����˿��̶�h�+� ���O�~/f�?WO���k�EW�_p�,�g�gD�2���5�������;�N��5n���g� h=d��-%<�f�`P�)��8K��Բ�j8��~�9+�7�%�������r�T����{�"�	� ��SHBK��ѨK��xN6v󴭊���Ju��C_�d���-��R�4��Yg����tsl�ֽ�;X�-)_��ߌ�
=�`���cl���:~��H�D&eݟ'3Tg��5=K����)؇�}t!?�����s��^�6~���g�����NU��J8�VC�Iz=���[����w����jx��uՋ�d/y>Ho��yVs,9���^8�|��L3�ڨ|�.�D�)���E��|e`�-T�U�"���jVa���(�$���!!�&Ju~}+��t�Bku(�(5�{��=[ġ�렢��bND�tf]}��a*g�;n�������%���y�05-D$#1DE*]k�̙�f�I�jY@�P]I$	�b��!�zuo-TyB#n��xf�gA+�YY�T�Ї�m`y���3><|&8��=��v��9�r@�i�lg:��iW��ٓ,��%ka�f�}yWfnr�S@4�U;�h?���=�׎�8��$ք�"#9IN	M�c��m5�����/�<�0��<g�=1��Q��H�62-�D 6��(AK��3+8�!j���.:5�s\�r�MA���q�B��jI��P�w�6������Z��j2I�V���R?�bz /��*��b�r��_Im����q=e�I��p�.�����_��&�#kBV�˄I;�K�]�S���t�O�����eg�#�$xNly�������:y�h��s<�e=-��qu�6��c�F2��4=�X���̏�L�DE�|�ꤳ3lM]�(Xf<���͜}�ED������w���]�_� ���V��X'4D�%��s�n��s���k����f}~,AՉ�`-�)UK�}���G�ܨ�\�?$����x�Y\�-��PJ܇i���9f]��өJ�lt�_WE\J#��/��V�Ց�2,��)<!�S.�� �bK]w�:�	X�0B�y>��EAd=�M=�.t�>��f�b��N�0�x��U�Ź��+{uF��+?r�UBM�A�#�:h�.�i3�kBbAԉ�����u�o�n*��m�xڪ��<���U�l��P;K���+#H=5�A��N�{�,�\�1�ga��l�9�F�Q�
)0��1�m#~|V9�o8���gPYM�>��O��� ����"ϕ�q�m�Qf���^�AA{�5�`�A�l����Lj�n6�!�g�\�i�2lw���6��;�#�����,��(������R��x�7�n��;4bH�y�t� $�Ϥ�탊�@�ࢋ�&���ګU8R��cg/,��sKSDn��� �I�����Wʩ���a�&̿���x]q�y�:nckV���a]��R�]쌠	&����t�C墱�}/�i����)�w�BT^�6�zT�jB�D�~t�2�x0!�m�Ej$b0��� ͠�G���N)�W��ū�L��No��-����
����rF>lF_ 
�5��	�j���g�s�J� ��dD�&,\z9�g�����+lMLRU#���i��{+���`*8�'���T�$�d������рqTg�*_Dy���j�A@wg�3�gJ��K�����2��pC�G�7��k�ϟI�x2�&�Ss� ����D�f�<��t%��(����
���t�WN�N��h���ϸ�
6&h��f�r	*�bmN"�\h}�Uc�q��~:	��4ҹ,J�;��Xv
����9V �jB�8s��\��+�R�vC�h�,!$�O���',=Êj���be�c���|J��p��1rn��kH��I�ς�O���e���${)�La_ؚ��!�虰��e�}��#?P',�JmHk`��!	�C�6��;ϐiy�'|j"7�ki��9�*��|���|�A�4�����Y�__��(���Ah�O�m�����C��D�"��Tk �½�}i���Җ�Wy�Gw�1C�$�&%�t�F��c���F	Cr����`�v����ߚȏu�Q�J�J���k��?W��"��nD���3i2*	�
&�w]PlV&6h/�Z����΀k{�)������?W����4�ۗ`�{P��J����-�Ĕ  �T�`,0]�nk���,�[.����A�^��kH`���#�V3N������s@o��N*I�۳?7=D��G���}��~�@�'���_�g�B&O.��Ќ�+�J��>�W��e	�-z�j�"�8��a�*g43�PI�_ �p��$,$����u�u��_휖���D��m+������YٱG�EI���ǌ����f�@ߊA�KQ�$��Sɯ�Զ۫�`_�;��P�(�Y��k@7R+ �Y�����ѽ�����my�U��ˠ�L�N�5�Ť5��}Ui^.Yo(��H�+2�B~9�\�A�V�h=u㽬*an<�⟱{�'"��~[�]?u���6�O�,)B��F�C�~��jS����5Dq ;>��TMn�����Wp��Q���LV{�V���S]z�Ӓ�sK�� @3CtJWG�k�&��Lo�?�v�� ��b��?����t�So�6F͒�������	[�L�x�����[XJ�'�z�� ֐oI��^��j��#����'��r��ǎ�'-�ZrJz�:֧��v�D������2��� ɖ�H���'������b�S�G]i^�Gq�2�����!�B�N�_k$W�j��p�?%[�S]x7D"^(�7�|����Y�$o�i/Ë=�������E�n��<�J�@7�;��r��%rC�\TW)�QN��+��S�8�'��/1�t͑߱�"��=m3vX�3A$6;Ra5�d�����6�2�Dn���;3d]k�6����������I�`I���Uu�[�[�=��Խ�g5fowL��|}�����G�fN�����NPn �a��7���*�! �,}#���tB�7S�6
���c�GǆG���
j#58+�M��Q3��&�wݕ�6��IU��*À���tk�(���?wN|KG����ћ�E��
*����.����
U�q��&VAV�ƒF[����G�}��O�Y���~N�����c�9(e��_�N���V�]Т
���\o ;`��1�Ԥ���ܕ���Q���iL������I1��"�؇���L��w��*��Ƌo_s\_9B��Nl�i�R�#���Z�pbT��t��N���ghk��&⠰9���
i�bo8a7>��p���B'��L�v��;�N�Q�C۫����2���]��į�����D��}�ӒO ���<;j8����I��SGv�G����W�sZ���<3f�뺦�"[��#�acEq�4Ȁ
8=�.�w��d�S���:��b~���:����'P� nБ}��R)(� @o�`LϏxr��tܴ���C5́�QیF�_|�D�"ǋ?�rV�
�w�=K��n��ݍ�P>��>D�X�^���o�J�:��p�]�Ėi���
�q��b�e�.B���ro��:8��B��w?A&N�~�S�D��;��)�i$Vϑ���N���K3"s���>��G�7#����y��~ܲ�b�ŝ��a˞�Y���ޙ>I�����%�Z���tt���X�@��vWr�B
��XpO!b��J�4Dg�#�wx���U�����a�&���Lŕ��P��^�J�(h���@���'�׌*ڼK'Ld����~��!�TT�Ɇ���f�*�M���P�K�|9}v ��|�]'�5�0en�Yb.0��ʍ[T��v�b6���L���	u�N�zJ:�O�t����>8�pيVb���.��1fO�?&_`ie����S}����H�WX�N��쭼Y�#T���u>g���%��a���M�-`��t��L���B�7PT���!
�t~�r��޻	�9�
�'�m�k�sg˱T���3Gw�j�l�Q�&1n�KL�)Bcƺ;6���֠?�8��U���G6�*}��&�i�yQaY���HVv��T �H,��Y]��T��}�	�&c~�W�ߨ)<��gd|;/���!m��Ӵ� �"�)k��o���k�(5�kH���$I�K���> ��_�>�!9pvi}T�����zS�: �+%����~
�8ܺU�N�0qG�-����C��"k���X,�����͠U�O�5A͛�Ɩd�=thl�l9왕��;��_��W=�)Q�,ɍ�ݲ��QJ�D�i��v5mh,K�|~�[& �D!~(��т$K�D���I�lcc'zs����_h�V�`�.hMoB����qkS���z�'�`���'����S�Uт��F����,�y~�l���;��2;`#����*@&���7�o�����逾>(��Ė��0#
�29�<�A���k��N=^�-LJ͂����J��yL�0� ��sRm0�Ӻ^ED<�L�ǈ���X�R�c��7�e����ܞ�9��Q/���=���e�p*�G6-Vv⤳S�t��M���'�&��R�C)J�Z<7�?�Eb�EI���Ȉ��բ^X1���H�L*�B��o��>�i�B4��A�6"x�[,�G��!󢡋WC� � G����F�ہzŭ�G fRGK.y�&ILњ&��u�(DZB��j׊��H�L5HW���\~�;�o�vy(i)f+�	�/^��]�t��H���O�J�$20���I�伞���X*J�qF�]@�͝mR�w\T�V$���TD�u`���p�|S�~�$sVD��)��QZ_���?.]6҂�Ǧ�����C�,�MI��)��>&����zh�W[���E�v-�����e. �y�ω�)�������.r��r���2�@�'��-Zz��?���M�d"��Y4F��f�_�ɌwZ�Jl�j$��@{���=��让:�*x.��
�z7�y�i�`rE� ��D�($��'�ț����-,x�P[�1���ߛ�}��zH��A�A0���%}����s���{+�y��"4��Y�$q�^cp�e35���D�nW�<�鑝���������g{��Y���'�ޛWZc��*FQ����'(��N�rW��FL�g�1�t	k�b"��ص�3؁Z�Y9��S�r��������p�g����lq��X�+΀Ϙ��u���{�mo,�C���f�����(�^���i�-�B9V�D�x)7��Ĕ!��8ވ��95%�5�c)���Mǒ��V3'�/�Zp��[�3��\�%�`�':_�#G+��N���q�@0#�r�C\�c#��-T暏,6�՜8�EL�a�ƦO��X7`�v�����l�c��������lqݻ��K�i�Nx�=�D���`�~**���a��w�~�%Ӣ)�]�,������ҙ��ӏp��6�B��)é ��-��2�bIHl�}�~��z��pPLå��I��>�@��~ŨWw��\�����Y����C�%���j�Xp,�s���B8D5ٚ�����O��"�"��Ҧ|i��0`#��]�`g��N�VlS��w����&�Qo����C_�W��;��"ΦװJ]�a�J`!�mXғ���إ��V|c��މ���C7SNN2�p�풁n
��f��Kƅ^�>yg����p�
���?ȶ�s�7������^�JM���V�24����5���&R^\;��!{�a�܊��TS���y8�х��$����B��/wis�3��1D#L�{��A�}��o�F���iFtY���'�a����e,�e�yjm�W`����ʮ%��o�zJ����7�a`��?�P�6�S{�8||��[�^D��ҕ���x��(NV�mB�;����[~"����ۀ��8!/:�v����4��'���tVn�>�k3���<��y&,��pJJ]��@���$���$�Bx��-�����{GR��I�y��dJهn���k񯝨C��%pri����5� 6�r�nP%��,��(Q'��
��)dv�Bv |9��,a\��Ćq�Ղ��=���u��.%�𿃌��x̂�	R?u��g�a�`����'� �WHA�� ��/�O.?ɬ^��\@|�qOFbJ]V�	�e��m�B�ʕ0B�^}����8ڧN@�Yl�q�ݧ<0�|��bCfB6��?�-�7I��BC�s�7X�߻�'b6���A7��}WEn�x��БJs�`3��tx���_�x,;�-w8G"���D����y0n�
9�&��c�i*���4��q\��m�DgA	���'j.�yZἝn̵H2�37��M��?��U�.���:�/bK*��rI^`��;m�9sj����=��<�SQ�C�^Q��n����JK�