XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Q8_3�ϴ��F����X��׃��D���Ii1	�ۉJ薥\�(\Z�����JZ����jRi��7!Q�&��E�gH����:֞� &�h�����7:z//��uj����qW�MN|*��A%���ӹ^���p�����gB�<c+pY���[�k����,�w`'�~��  =�]j�q�ޕGWASU���T{���@2�|ݩB�2�k�I(�`�*�|?+ClQGo<�����݃ڜ�V��0�T҉mˊ�
�4O�r��U6׶<˟�T�L����̨�"'��up�*i4�o��b�a�e\ͩ�\A�`����[����p*��������cd�W��vw��m`���Ƶgl(�5��g����MK��Ҁ́`1�E���?E��K/1���yp�L�v�����-���x�#CK�0]�V�I�@IW!�Ta/�S�4׾fم!E��6W|�^�7*�@��k t娠)�߹X�C�ꓰ�%r���<�`�@��hׁi}NϽ�8�8��O��[.����~�Ƃi� ��~��Q��jv�^G>���	G�ؕ������#LqmON�gI���L'�]�Ez��󗟓��O[JR^y+3'��	���������d��X��c��(�G4���tɩ]^��n�Y�
��Ֆ��-h�,V� W�� 8�AiR�a�E查l��r�|?�S���ify�
�<��U�+ ��?�Bv�J�	M�,[�.�w�	��j��cԨ�����8]XlxVHYEB    9efe    1be0�d{�`�1=B�8.�exqê���u(=:�]mO��`>���fA¯�L�9�LP�� MDz�Q����	2�Uԇ�`=��߾
�v��4ᔰ�$��F��"�9O
f�p2l�Vjt���#�~_�w����=��V���e�K�DG[Wk-�;^4�n�lx)�q�N��&7�j{V�JҲ�WCd�8�*�1{o�N?((�O�8��쬅�)�o|��>��c<�uS�Vw|�= V�_S3�)�$aܣ�Ef2�4~F|�Em$.�R�aN�>j(=W�Ŕ dE:W{�vMZ���P蘲T�����������
?��lJԘ�*3�C�d9$���^;��l���?��dۅ/�H�D��o5�����G�0=r#��ϓybex�rR<wq!�u�WrR#�����dʒ6�0�Ol������@��@�u%������1*)�M��5�%�pQ�3y�d�;+��(�[սK��s����,+��r�pE�n�8RnO�vt��B��JY��9��u���J��ؕ ��kr�ѕ3�c�q����D���xoRO�g�^��Ǆ�v��E�<�d:P0R݌��⏐��~4��>6 �*��s��=�6��!w�QR��ѩ�2|j���1�ic�H�ѫ��g�1q���˩򰤕=D���<\�ᒯjy"�Ģ�%���/]��cK0��D�+\BA�l̖)2H�(�ۈ���#�/jk�'s�Lv[2BCCw�\�>;��v	��(�M�jP�i����K�SlK���p�U���b'�2�FnS�zxXp�
��y��7�5N��ٍ�S��(/y.-�TvH�9+\�V^-'OU�p����}>��Puey��DȍRR�۫vm�
������:u����T�%F[Ō�r(����|	����ޜ�n���	y;�S)�b1P=T��G���_��~�.,G�qbe�/�/
�['���/������+%H�]�垗�]�Zwg�bz��!GbK�9�X���|��e��D�]�B*+?4�[n���9졡���	���݆���}do=r\�5TĄ(�{488���ǓQ9��ң��8�����˚��TS;��1����u/7F7�3g3��̆�pR�Xθv	�rd;����#�	#b�5���3-�;��B~l6	΅	�PuC��g}
��4GP'�!9�O�Չ�	~r!3�Z ��<��1�{�D�����K�lQ�]���T`SQ�,�S�b��yc�F���׾��r�?߽�S��NfRt�%sN
	D�n&5k�I��X��ߪ�L�#|'+��4��M�A�V���=�Z4zМv	�{"#P��'U���6�.d�b�f����xΙ�OVh{��.�kf�ܡ�/�Ba��L��a͉��Ō̚��*5��N�'�C��W���iv�ѫ�@:;��w��Ɂ+ fO����!��	����u�D�'�duc������8�w-4�L�����U�</�>r�Kfř�4ǔd�i��bV�OE��r�;��$��ӌ��=VH��٨P.����ц��?�%�����t��]���������4�ډwL���
?7+��9aQA���bl{��9KV4C=/E�c�N`B�]8����m-Y�B�?�+Tq���c"� �S����	����Z[�mT��Ld�{ra���O[��P�dC������Q��!���ڒ^��¡;���ˣ�Բ�kP�6g�����>S֖���91�1������q"�z2�����]���mZs�%5�j0(�W@� ��;���T�&(ʾ&����3��&���	'���5o��h���+�g40J�MIy���o@��X�V@�)/l9� Y���}A
�V+>��N��}���h��h���p��dE����uh�D]A���MK�uFT�Ԗ�U*��� /`��b,��C�磉@)$!1�؜�A�I����g�km���ߚB��𱦹P����ڙ�]��-h��]��:91���^X�4���eXHb�FT/6һ}>�-�rd���?�=�r+xxdʅ*�hW��=(b��/-0��M��I&��ٲ��,#vD��S�@MR:g���m��� h���z�hN�z�Y�s{c�8q���H%ߺ��|r%x�;���ć���_���X�>Y@0�}��S��,��ev\�:�X*�0]���F��̶A�4�2����� �P;	�ҵO{F\C�4��/���U���Y�;c���ʃgU~��`�X�gc�o(��'�}4̉�sH�I���7$���W���f��[{K��e��;hD���&���8�]���[R
8��
�_Q�wq��r�������e������-��J�ɟ��g�.�!��m�X��_[^|#�M.�>���K�6�S�E�7�FzK+@UR�R����2�c���htF���,��B�XP�d��rX���hX~M������WF+b�c�C�~�1> ��-�P�1�f��İ-{N�9yJ�����x���-\�z�Ԏ����B��9⾲��I-g ��ֳěA�dH��h�������v��%�T��a��NB% �|�Hp���k9]*C��^YCB��x�D�F�!���.�?o)i4T���W!�l�d�0����W�b�N�#-P�?+�r�����>RAx>�T���EM�@5vDEXЀ>j�n���d/�x��]=��.��m��'�?��0�h��_�>p�n1+�+K�6��x\տ��_WQB��xr����ʂ8�~s���v�QC��	h��`#��Q.�m
�P�v��~���b-51�M�>g;%h�\'&Rl����N�&�&�HQRn���!S�0�fK�&�):�+�)�w�Siy����`���Y���OPԋ�LW�T%�fJ҃�vC��J�.R������=�픪6^��o��*Q<T1�t��?k���Ǟ��j��"�@,`��6V>�E�-�G��+U���v/A�˃�����ňs�@�W��6�*[
�o���oW3�D���؇r��ߵ�{8e����`�Ka"i`�h,6�J@���}\����G	n�X���!���%�i����J�K/�J&�׌ȇ����V���T�����ݴip{c����I+D�� s���]XV�Y8��5���^�	�5���[	FOl \�HTi��
�z7�`ME���k��k�)�ʻ&wʜ2M�UH�j�_��^,<Y������u8���OAi�������8�&+J>�1g�Ŵ�����y@<Z�F�.r�ü�Z\�'s���+i��mg�W$����jށ�w���D��D��&?�Y���7�3�D���;��=:,n\����Usj��@u�#B��Y��T�C��UL\{�.D�4����T��^�j*,h�H.Z��?7aO��,�.��@~<	o{k.�ɝ�P���j� �%�b��؝^�0�<�f��%T�=t�E��}\Aϩ|�^|��$űF½�P�a���,�,�st�uOA��B���1|b�8��g]�N�+�@�k�%Ue���?�0,0+�G��;-���窓�es&����3��5�}��Ӓ�Xz�8P�G+���#:_��b�_�X7;	1���u��@ì�eXZW�@U�eb����|���a)��a�����Ǎ�t���W[>���x�ɮ�2@>��X�Sh��X2�V�nk����Hעo0�ZM�.�S�ߺ2��d��_~Ҋ��Z�N����kadX����<���ˢ #�wl�+ӳ�!�1�k�iۚ�Ѩ!��;ڰ����OԨ�.�ui�s�d`k��t��0������\�X2����8���ć�>KoT�hnbO����Ǜ��1L���`��$�z�����U�@���K���W�~��{�F�(Sh�N��j�$�>�&ҕM���F�%�@�Y�P�/2~��:�男�.���L���[ԂѮ2]�*;���Q�گ������GDo�}p��`�!�%
�`�y(���TB�#n�˕��w:\��P�!����a3d\����{��+���Q��1 K��&u+��·��J����DxmE1��"��l"Z��F�d� z��o.2͑��ڃ�3X�Xx�z׉(��@9��[�DiD��W��Ʃ�}CF�?R��ǈ׃�����:H�N�B$??�j�*�j0�M���BL!$I�t�pk��J湰��^(cc�7�I�7�M�
���͛�����m8�찟�ET8�����?I%�+9Y�zi�8�XO���h
���Y?�/��� �7t�Rc������y��c�Wk~�ت�D�Kr�FM���)��|c{U��*�6}�Q��`��7g 淴��1��~M
�Qܘݽ)V���N�K�H�*}�K�f�z i�G:�$Y�L��˫��so���2���nkKTH G�2�T�x���G,�P"�ec��j�;���/�7�#dYy=@%8{v�a`����4�O���88�7���*
V����DŶe�z�Gg��i��{�-�I��x?��R���`�C�v�����-	��J���{�L� ���D�YІ��zD:)R�C=i3�+�ރ��R95�}J١�!�F��P�����8�o�E}�r?Kz�SA�������Pj���F�pC������}�j/�.[��W6�,2�QX6ظ)�����n�9wKB��_Ц��p��)��a�]��^�ѕ�˻�F!'�+���	ƌ������GBz9�����[�q|���w�'6�H���w��C���Y�"a�X^7�Q1K&-������p]�R갗2�0үY]��c�����*e�dgV���,VX��~�t��FBl����L>�L�Ð�(iBy)���OY�vZ9PP{�#/nD�33Un��Vs]b���� ^v�u�h�־^�(�)!���˄�j�|������dֱ-�I���H/��Fy#��/:�j��"���f/s���X���~�d+�9�لH{s�C�ү�"pD�{c�7 ��sꋞ��s���=�W.�;'<�ϋk�tk���9Y�WKlΦ�$���g#�������(��y佒;T}�U�{���g��S���8���|nv9H�%Y����;��bq>�L#zT>(?�
"!�6c�w1jq/a���0r�b.d٥a[W�4j��L���<�p!H��\��c��ӯ���"���x>��,g:�+E��&2�'�������.��Wp�ż��ɝW��h��5k���,*J@�ͬ���2�v=�	�b�o�>��<��L�R,=i��W�1�b�)�>'�ti���!~�̙!�b��q���u�*#�L����t�RlO(w�GHHU�9š�Fݙ$Xw�^�Kn��~3혆ޔ�}nn�V��*de��}~\A��ک�r���wSS�9�e�4�ܸ���Cp�!/�۞�M�j�J#�7��q����^� �ӵ�V9���4��^�gۘ�3��Cy��8n�Pro�n���.efHc�W
Sx�?�
ߓJ�J�BL<5_�=�sr�HaaN�P@PT8�ٸ�mE%&�c�x�|�3���M��E�)@D����,��K�v|=��{��j�C�{~C8�,���B*l�e���Mg�����9j�eo�+��q�S��D6��|:���7xP� )�3	)P�,Rz�K����şBF]���NpĖ�ʙZS��ֈ{8�G�a2W�-�\1aX�� �Ɍ`p�Z��ȭ��$��ԣ�EA*��pM'5X�Nɹ4�w�\���悒S�P̕�I�=������J	�>7!j��u, ��=�BU� !Ծ���6��ǷLw�=R�Xm�H%AY��oF�1{�;ߦg�Yաk+�e��=':����+��I�^��NKč6�N���M�jތ��pn
�m��v*�o�ߙK�R��,�V0���?��	w�_掝h�2�~���`__�aܒ���8��slm�%�i��	D"�����D�p2��P��l�!\�Y
��� �,
@s�?��ׂn�F֧�nXSXiA�lAf�f/���J(�����C����;���q1�6˹�}ͤ�O���N�ߪ�6+�rFL��c���0|5���B>�~��0P,g�� �LC��-!?S�Z*Ϥ�"�tZ����V�f�A�;BaG^IP��5e����7�?|`��K��X }d�C�/B�4)�b��$iOX�>pf8`�ie�5xK��r��6�A�����{5@uԋ���ۆ2�G��I�����=���&RW��;r_B����=��*^��9����']�B6��� �D.f����")�g��`WQ�ɗ;�Ղ��'n���M����1� W�֩�S�å‪"s8�0��M�����yhe�n�qUU��g��4r����Cx�>�%��C�	:��?���UL>���'0�-��#�I ʰ���%������.F�$t������9L���Re�k柴�aY��aOH�6m�6�=O�J1ķ���	���h@�ƾ��$u��>n��2�(
0QX,?�槂X��JRu�z��+I@oA*ǬM?8�I�q��S���8�N�7���br/�,:~��<8ϔ롫�6�r۟�l���3
�`�� ���pd�l^v_�5#�ɐ|����J$�(X@��&`C]:�F��������L��Z"�y���J܅�T�H���v>�C�?��#t��h���	(���4qgdk�1JKf#g.����X3��c(��޲{�X5c<���(p196�0�/,��
-`�FLI�#s**zoi���p{�_gb��4|bW,��������zeS��Jb�q��f�6���6&#�i���&D\ڭ�a}�*t9�>a=*�9W�)H;�ߐV9xY��y,tC,�(�3� 7��q̃���f�|oq�Y�5��p4N������c�������+���9����`��]�O�I����?���A��B�	ر�J�i����j?N����\�h�G�0�ݙ