XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����@B&m�h�5���5��ڥ���w���t1���v�{�'7d}����<ub��Gѓ�}�K��jV�r�7�Î�#t%]�<�)��G�yN/�Pɧv�9�b�Q��#�F�{K�1>~��X��@{�ѿ�a7`���Vu齙�E��Q�;̲��f*쫻U�=�ٯ�3�R�KT��wJ�"����?��T�-i���0�g���C���/)l��LY\	�J�R�Z��RiǕ��ʏ�[����6�>ma �́G���b.;�"ݥKE�����B��$n�L�0��Wp+�ѦE��¬�99�
kgU�Tx�'Ӗ�"�b������P/��vy�+�9��5�K&/�`�Yϑ��<����N:ݯ�>^.��}����G;(���3뗭�'/O%��+QɈ�r�e��G��l�|�<��	a��rP)�μ���|�\SrDSћ)N�RQW�KG�q���<�)�#�ą�<�s,�&d��5{��"�$NY	B}��,f����*�=f+J,�|�s��V�5D����ܼ��6�m3j��/����f��DX�f*ɍ��{gr~�U(,��/��5�U��{CLެeƊ�`ֈ'�V���WC�j�z��!=D��[�y0R͕,);%���c)>A��N3������Yi�z�]�N����A��"'	���.vũF��	�@����R�i����;�lFZ㝞�\�Q��,yv�-٥(��p ��`��b1S��Y�p����Ǵ)i�t}�XlxVHYEB    7187    10d0�g(��x��ի�,�7ϖS�o�Zׂ/���{�(6�k��#���6Y����b㮲�ǿп\
�*��)_�Sg�J�����l����Y�lw�� y�l��ŏ�y?Dۢ/��|;�aꛩӱ?�Y�կ�R��4�QH�J}�DR��zV�p�o!�z�e��7>�&~�>ҩ�k�?D�4�����O��������~@�%]����v����j��QP�:Aw(*���v`�5o�?%�N���03�7V� Ȥ���F��t��-�5�d��T�c<�0*��}��[/%�?=TG�x�7yJ�	꽴�'aJ&u��f��8�o�#���m֕R���&����8�*���2"u�7(�B~������#�j�����IXܩs��0�Z{.-�OJA�]�C1w'Ǵ��B��d�#��4{q���7x���h���"��!�7Z3�S�cc Z�{O�.፳����5%;w�?32e�c
��9s{\4��6� �h��c��b@drЀ�eP!�u�T���3O��{����oG������YCi\�z^���t/��.شW��Tv\$�bٻo�'�W�C��J���Uj2�ީ��b�[�?�hW��!vGx_O$���J�7.�M/f��A�1��Jp1V��F��R4��f��)g9`��DA��6P�A�2(kK)���9R�	���>�����]+6��m>l74�BMUG^���M�P�'[iƥ�-�@�w�x�A��q�o�w�s���p��O�Șl�O��,���4*-�6���A�����BRebg�BDi��!2]�k���S^!D P+K�i�� ���b[��`�L
�)�Py���,�l���$h_Yw�&�WC����
L"��Ͻ;�&�6�#B7&��@��Y��_r��t@	��W*�۬����y,�|�Qҟ��n0�,h��-��W	�	�*`R�_(��u+�P��c��FZp?���ٳ6G��u*ls��QN�����G�T���3�A=��p��}���͕�HT��`���{[�����y��e5G۶{s$(�.wvupd�4ߕM`�r�F%�y� [������\!���ZM�BR���W��i��᱄�og�����P({���Х��q��:�
S*m	���:	9O-�5�:x:�즿3���F�Ѥ<d J!L$��(��PH��vͯة@����&Id!$ÓaXTG{�PL�qr+{�B�9��YG����_����5�	���Q�Z����F�A�����@�Ǔb�'&+�81OGu,T*���fg�<��d$H!�:XV�Mpd�3�]"0�ʴ�s�l��$_�f�D~y��������!qv}U�1�r��7V�� �NQ-c��f^e۱��x���8��|;�ճ�8�~�!?� �B�1������6)�a ��[2��5�ޝ�_�I�]�;��4K�'�h�Rv[��0�KIARv1����vB��]l�`�\c0Y4��#_
hk<��6�F���<?:�I����q����;�Y���)�|�t܊�
�|u��`���Œh��|���2D� ����ܷ���G��'����?f���B���z`�m �6��u?�v���:����g`�U^L��K������B���pV���V^d��c9"�Ή!����A�ȃt�l��E��+&�%�#��9��������[��c���g��U/�$*���m(�W�n�z��-��6:�r�wwz6��0٬�HC7�ɺsVsIP��uMs���]s�$q��N�*V��U�7������H/��m߿�+�H9�����v� ��A�0#X5��8"���0(S
��q��?�\ȴ�#	yI�W�ߊbB�m2M�W����!����Ak�±�?���;F�Y0�N��UfK��L$���#U/�q�x�>}@:^=��IAt�efvb������!I�GPrK��5�h|���(x�	�"�eu�N�z,����,d��l��`P����ad�L��*`�wjWRt�љ�C=��9͌�"�����:פM�;�􇩫`K�m�<׏�"���9ţ+�r����ԧ�;˱=��t�ܹ�f��u�+vQ����}O�q�C&<��P&�[�K!��h�LC��/�rP�~��LD_�W������ɐ��F�1ˌ�g����[����n�4�v Lg4�X�H.�V���p�g��4_�1�-:Wm�	Y"��Jvvk@�-µ���i�=���y��2,\�������/�
�6��崘���U\�%`��hƹ�(���������N�}y"S:�5鷨ZB�w�MS(��u@�O
ƹ������ɹ<M1��R1 ⢃�}S��Ea�����z+�7�g������/�dTAh�˧\��5/�m �ZS�[�t_�D�4DN�oE���u�x��/�Mp�3�X,M�����4�+�^y��2¸��A�|x�5�^�eH�DJh�L�@��\�ɩVl,YT�͞��hb�!�SQR\/��<��zsb�#�?p���>o����U���N�էۺHDۃ�h	���@��a�$Y2ŧ^C�]�^HE�e #�=JHug�z�Y&����[������ɾE{ǁ�?bd$�%i���]<$�QP;�Hy��~F����w�i��$f�bx�t�ZS&zZb�h���f��b�ł#���gO��W���T@�> ����a�f�n�/�qI.c�g|8���j��M�����s�����Iv�bZ��cm8��}=��3j����K�DT.=�<b�ho���_� q�Y�q<O�ײ��Н�HO+g ��`5�xH4}�O��o�]�e&7ݳ��H+�����W�����4��	�l�_���}�	b+�606t a���:�n�ѽ��~I4N�~ُ���0��'DxB��{2���:�����H|���er
-�YnZ�(����*OX����\:��{�'�{̾��d���~��&orА�,�nk��ts�(���V*�HM��޼߆�]OA�Q$���P��c��uI�b����g��1�r��5*0�=k�ow͆T8}�:��.�g��PͤyDc�'�'�%;"���`�%2ܻS���pH����G�I�a�Bӳ��gL�P"�c�h.ҹ�PQ�cs��,f�Z��˾��/>0�W�$: �X����K(�4V�z\�T�����¼�]�dp��n3�yFs�LM���՜zF�Iy�ρ�ɓ�n����yvg���J�U����]sܹ��gy4ći$XA��ߏ3�N�_����Qύt�)N����OD5$�72��/�f��1���6�#H�_d��8��ڋ���]��%[�I���Y�5���J ������?����I���u9��%EeHR7ߡ+O�;VK��S�3���� �kZKy����)T/�Ic��: O���K��[A�+���#� �� �6��$�acL�c��3s��H��
f�p�̵�����O?�-�z�,ODh]���}�6?ފ�jO^xNkNJH�q����nvc/W�'o?�$���q���
�R����X���wQ�xs�P�m��.�~ |:?��2M�
 W���y&3�ݛY;�햕3x }~�!b˻;f�q��^U�܁9s3���gC��Fm?f{�-�7�6�e�	�K ����zuE�a1j\��Cw>8�L�|cʾ���G^v�Xhb ������o�w��&�x��iP,m�Wo��.�Вd��F{,y�/��:��iA�K��Σ{>,��2��.�[O�|f��Z'�����t�����e����Ŋ8���":�[�2k�� �DIی�S;�`=b��'�E�������,R|8���v���M�CK�(�[���֋�o�c�,��e�9�����-0O�e�'E��)'��I~3��G��4�Iц���������֍��f3̰K�sl�I��D��Qg��>���YV��Jn��Ak����+�o=��!M��1�k:�P%�?=qAkM��,emT�Hm��+٘I�;�=͡?蔛؇�B�����&�dP]r�e�$��b��|}�ck�@vN)!�4���s���!���/�[>�2���v�cK��s�>`��5��B?����
�*����s&��\��o��"������_���Z�"��Q�J���K�Y$�[.�M�y��f����.,��Py�м&��-J�s��|��((Ʀ�ֳ���ƀ�f�7�,