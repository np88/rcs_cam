XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��3|k�ҟ ��K��������!|5�`Ո�`)���`ȟ�c���{���>ʬ�V������*�p�8��g���&#�+p+X-�5B`-~t1���4��a
`��[ q�D�D�=U�@o�Pr$D���.e����o�?x���IP_~Ua����ea�$	��ס����O3��F���9뗖%���H�����x�X�gzWT�狖]�):w��|^,��}�jo~%a#rX9Q ^i1�x�X��:C^�+�+`Q����lm-}�S������Fa$M�dA�Q*�:T�r��`Hmj�o�r2i��R��f���-�l'J�ճ�[��o�V�����i�6��VGx���?ﯹ<�9�FG҃�闤���ҽ���g�w`Ck@����oD����c}��j�/��Y����[F�32^�}(X��s�
<0\��k�������u��1�pNM����$�-d`1P��u��^d���Py��
5�ֽ�xB��Z��e�J�ǐ#f�C
�*�!���u7�R����2'��JD�#AH�L���h����*?ҏDۦ��),(N��������w�~x�6H��z��~�Ѹ���ϵU�+����e^��@�����u^G�*��+5}z�s��x^k��]�v�q�3�P8�	��n4mX?4}I�2M�.j9��%[�e$3� 8��ry�_'��y�Cͫt?���zd���;�7��5���M`]�7�ܱ��$	��˄&��)KM�0���7iXlxVHYEB    fa00    1ca0���_�7�@vV���G�0�X��61����	�����ؿ����?ԧ�`�ˬ/��X�9���Q�I^)-�׀��S��d�.bB� ��5���e�A%m�X�ZRT��m��J}�l�D�gK�~	/t
����W�Ԝ5�����n�Qɣ��yB_��Fy���S��<�R�\���#C��6^4K��~�m\��L��g�����+=�z��\T}y��I����|��%�>
�D4`@�q�(O��\Y>0Cg����d�����䄡�^��T�X9��֣���Y�;mjx:X�! @d�9pq%� ����1����l��*x���؝t�)?V�]��0�ȕ!`�z���vߴ�1F9F���63f�@w�q���5�F�N�m�}�o�:�SCs��ɚJU�p���jC�W�>q�av:Zt&���W�ffU#�������Gk��PhR�dp���|�!�('��t�ӺJ"��=�㴚qf�x���G�8k�[�]9��5�0�v0�,Ҡ�B�����1�L���FbE���MH2�A�>�]�9�Aq��0{��ĺ�����+�AD�y{s5�[97vHkR��D���,A�;��?}�#y�e�y��� �{�A~�>+#b낆fH��㲱a7M��MՐ�d��̇i�q�CŌ�����l�
�X���Wr4&�S��A:s<L���6=>���,\�]Uc�xsȲ7��b�r(�����.EK�bD.Ԇ��Cma�T�=��eA���:�6���r�F8�3[�l"��x���ߠ/ �zTB]u�Si�pob��n#uG�1t%��%�ǙҬR�19�nx*��3�U4Z^�`��}��O:�"^ၫ%٣�hWb��mK2�"r;�����qF�@����σ�y~�~��[ͽQ~_^��}�u�� pq��p����N�7	���\3���F��î��4>:�� �5 ���4^T�т��%�t�����Y����6{X�K _�K����R�j��e�o�{��[uو3{7eĊ����)�E�W�b�|�����*��/q2��c��[aY��)�b@�a;�%�q��iX9���3����� �_��-�1��q1&�oa�e.B�|&9����B����#����a��vYq`H���2��3.����I�I�X�`l�@Z7?���a�c�����;y�]�`C���*k�<���JZ��[��2��+}zQ��(_�+�yB�]lz���ō�!E��+��&�	�6��`�#8}p�S�7���;2�,�����P71�E��H��&���H��U�¬u�(NBa,�G_��t���3�0�s�qXO���\��I�j`|�B�߲�����l����o�@�GH6�mZQ����7x�XY���~��� ����f�u�������y�w��]AJ�u�Y���S��2��_O,֝�	`�6<��pKVH�\Ptt:��1Q9��}p&.�C����7�!>�-~e����SI��nY\(y��IT߸�Ν1�{J��!��1 �+�Z
���������ܘ�ȧ�B���l34�q�5�Al��H�d=H?���0`ƺ��q�ޛ���a�b�{C��=a��?�2�h�ɷͱ4���[�}�F�WbF����흠4���o�
h��a��#�YgN7���Ω�!pb1����#��g�e��n�ؚ5x_+m��j�~����,_�@�$F)�9��̵|�y~*�1�G���S �B@�ej���I�Y�}�a�ջ��Ѧr>��i���2Ѧ1����B�"��ͪ4�\	�[���C?�!�glbMa x��A��{?o�'��0��&�����k3@���d��?��$Ă4�?$u��tK;
2���&��S�R1���m�ЕQ/�Q;j��@;��kc���:k��k���tkV����]a��R�!�eɯ5�s��0�B#��E�*�6?m�Y�<K�,hWL�Z��2G�y�QB9�Ѥ˳�H�9�u�!���X��[xk���Wk�'��������j�H�Ml��(3��OO�H�2� �g>���D|�����je>�W(���W�������2ʛ[����M���5��H���B���ާ��� 0
p�,�P��ҹ�/���K���Ĳ��E�L}zV�r�H|�j��Ц��"���
�JV'~: C���b֎/)�̀���	�d.�� �g��]��|���í��'�V���?��1�p�S����	��(�N(I��D �g���4@�������<��O�ȹ*Y�ʚ�o��N�>h\|p$w9t-M��t]��Z:v����m�δ�-�2��(�a�}���w�V����f#�͞B<��i6�Yd��D�Ն�3�p��"�^K�n�o���m��͗��}'�φ�M�V���b�u�F@�A����?�'*�e8���~M��u�)ԗ߿l��;0�U�G��O�y>�Ŧ�$�nc~������J��L���z�oqJ�LMT�g}OO6���Kor��'~�����^i�.����>�a%���~*d_R�D}g���8�B�8'+�i�!�̣L�5�A�N�$�.��<F[�F'��p��y���
X�vL*� ��ٲE�\����(,�����ovo�y��1��N��8�w!S��+�����H^o�>��n��	� �6��F$�|ԝ���r0'J̈́?���y�R���H�pNu74���{ar�+<T�I�Ű��m�A~����T�~s#���-��-
KYm�@���nJ� �����z٪�<)��/?�n��k0����B�x�Ĕ�nP�Q~(�i�?&�̹�hӣo��9u@��BǙ��_ݗF�8�d��h�ֶ\!"��b�6'ҏ��ؚ4�k:�j�����Ҍ�)<�A(H1��d�!�?�����Xqp�#����=TR�I-��E3�k{��_گN�9;��u,>3�*p�
���1n/3�U��^�F�1�v��TK���i�7ΙQ��0�t�g������]~�+s����/���J��º������W6�g��eł�NN������wD�S����+�R	���u�������Biv�V|YH{'z��®��F{����k�"�:�*&�e��֪�u��e��N�?��y^��%����؍�	-Q��&���e���D�@�O~�3���G ��
�z%�OF=��@��a�f�c�i���RǶM�u*@�	�(q�!�e��d៯�]�����PFsVx��X���|���#Ƒi6iS��Vx֠Cb�.t�h������#1N���'f�I���!����I|4mݛFX���q�.��i�V�O�#̱q�����B#��[t3��m�vjӲ��Q�L�'�|"�q�'�c7:Ù�Jqݍ����6��kץ:�C�f������S����G�3� �ux���ޏ�M�6�u�z���#�_�u����XY����P�dd�Z�U��SS�xG<Uȟ�����~8g�0�q��B�>�Do-�������i��@���(�{�ߞ�xQ�����}���Ԯ���M!k�/��^?�Q��9���t��ä���.i9��h��,J��j��u��w�B؈f�Ǹ�/��/����.��Q��ݹ ��z�� ve��݄#O$wN�����A�;��;Nxt�}KA_P����.�vi~�w18�� ��0���8�˟��]d��74R�"����g+��,4�$�]Ξ+>'rG�Z�q�������W�� ��8D���3�T�#Z��z�S{�&�./z}�t��ixy����H��;8(����w2L��0�H�ƋHI������\�ɓ[96L�����iE�Ť�͏>ԕъ��O׈�z�K>ނ��=�nՁd���L?6���n<��G��J�4�3V�������+�G/zĿ`<o1�(ŉ�v�1Uu����A�k���/6�I���].Rd����YD�$�טYc)>$�pe
��	�OI���}�_�=fA��_��w���� b�k���&ER��6���]��S���nG�sp��nk�q����F�0g�0S���V G"h']��Z�jMuz{W1R���3���SN$ߞ��K��eQ��CD���'�	��w��m���e��0�[�Z�ӥ��1ireZ��=]w���#��A�w']���(������`[mG�e�����Q��xx���r�+3Jq]p�B�nd���Ζ��L5zpa?
��� n���sM�=Z>xzm,/I� �KO
�Lrb�)OTٳk��x�G�1�$�q���_�;��Ҫ�!���fV�݀S2�m�߶b�v, ��Geח���
�ق����i\P���%���C�E* �PL��:��Z!�W�嫏�T�c�C���5'�f�Q��D�#�Ŕ����J��9��F�e�ؙ/7Q�;��� ���S,��c�~�_�!V5�	���-Lk�a�vݶ!�T-:�x�⹰e\}C"�����1���f���(����)�	�v5�����@�ɟ�C뉸���bMWF�4xJ��i��}��ƪ�A "s�w�Hۂ)a�:����7�!:s@�f�~{P��V"o��H�ZB;�#6���['-#��kU�x�4� vӜ#��X�ؕ�4���DyL��?W� �Rwa;�h���0e��34u6A�#��X?F����v\�B�����L��9�`�XWw�_����F�ć�n[�~Ԭ?� ?*��g82��G�Id�w��b	�L��}���^sJ$6R8x������*)�o��t�@DB���XJD���S��n���j�J����N�O�gO��V�~#��SSm�]��<�H�ÈC�x��]��W�Q�	�S�;=U�{r�^J��t(x0lC��8+w
^;����Va�ϧv��Gy��g�D	,�֑�/np��Px��E��&�� ��k}Z5�>i"�s$����dL�	e�+.6�o�K+�ˠa>5����"���9�x�!Jmb|E��u�B6��a�gNr�"��<��;�Y��&�ј6)�ĦB�B��}��}v����E�.��W�r�S���+�ݘl�RN��W�c+�@�Ba��om���]������L�y>t������*yg��⥟����و>�&�xā0��ycw�_��J`>r����R����caJ�����>�����U�'�̾�J�}���$��0mA��#sm�7�,�b���,��,qu���d��-ǻz_�/�u�>��D}4*uQf&/�+Ŝ���,���6�A���^nZ��8�O��h��S�A2+J�fH�~�[C�F��PAX��+�3 ��Q+��C�%$���~Hamы8��]Oy�,!�J����ڣ->Χ
4xB�~�RD��w�τey�b>��W{�7���yBm������R׺�C�Vk'�V��Z�.�����~��'N*u=!�G�<A�|�,�(�e���d�=�v���e�a�X�Ȥ�϶$؝
�pG���Ǜ��	������=\�+ض�bZ��k�=f%y�/�`��B�*(͋���s�Ė\��!�
o�!�?���튙!J��,o�%ǥ�ͽ8i��I���odN��ɵy��Fh*�G?����n8�P B#��m�{�̇�W���p�A!��*�[�9dL����l��}6���,�'�'#8\�s]k�p��+����&����
B�[r\ml��ߠ�=��ɡ�~5����h�z�����1t��kϵ=� ���ֈYJ>k�d@!+&ɰސ[��R ��}=�6d[�ehՕe-��x��ڦ�?�EB=�t��2T�N8��RG8�{�|�UƳrn���/��q�� �ȃ�$^fM�+xp\���`n���/��1꾝B�*��i%:+�NS5/cXf�0���M�呌bVY{eq��u���ќ��X�g��!DX�E�(ض���_[�g�t�4��yY0�f��m__+��,� ������б�r�sE�F�Yj+k�z���y�υ��if'Ȼ��>M��.D��ܜL��W��?8?P�1���3���__ks|�����v��.پ]�#���0f�pG2X�f��D'�^�ɍ�� +H����ٻ��&���ݕʓ�ld�QSצ��������2���Ƙ�%u0'�̳�䖦Ȯ,��M��?��Fo�0+𵱕Ȏ���¨�Iq��HWJ=��es�uR!-�Xv\��+�ph�]e"��ē����N�r|�N�"$jQ~N��ۇږ�I�1{��b�Ugh�(�{�H�Mk����2?��H�Ę�/�exT�0��2I��<���s��U��p\����hH^m�+"C6��t(G){o��(hcñ��K-�oZR�t5�
<B�x���NZ+|�b�,r1.�J�ܶpY����9�m�o4�x��1(�,��9��UF�ᑛ�Jf@%E�h۠wPC����?���M�%Ѱr�9e���<v~I̙�J�&��?;�Z��p&�����|?7D{�=�=�J�_p�+�|�5c+v$�C�wҿb�|A�e������T�h� ��Z�@"�^����������ʨi��,�4;Hj�P�}�Qc�k��ԔE'���x4M�b���v%�%��m�@,S�Q��t
^�@����S�:���~׷��Biy��`�k������H.�pL\���׃WI�"���_��缝�
���^��'����sS;��Am�a���*7�������I��1#m�ڈ��?&{yQA�<Qڿ3���X B�ڨ��B�G� 1%�n�H�@./����9(�-A�0��x`��"���̲�Jp*�gB�������Ս��v﵊k���~q]Ӡ�R�6+#���#��[F�T������k�ɪ����k�*!��灟f��Ә�_��WK⌚�[B�]�e�f|1���[fɯ��Jt���gO��W4,6w��+ϻ��B�s�b�	��9�M���ܑR��W��Yc*��ό-��,i�@��oP����w�=#��4��N&�]	�e�Q(��iPc+Մ��դ��g�C��Z��~�xt(�������1<0_ۏ�U�(R1� *P�<�<nc	�E2���*�gZJS՞1�}8�Zct����gk�8I���EG�n"$ k����7�e�rKOl&*���I^`��"�Q �k�k��V��V��K�"@_�:��vXlxVHYEB    fa00     cf0j���I��S@Ho���Ӷ'0o�4+�]4["�g���"��$�Ì�p}����h}W�ӹy��&�e'��!\~ E��ci��Vg���	�W��Ϛ	qLu�H�̦��<�����iR�My�o�K���u�8cx�3�T�<E��~2~PY4��T��o����F�I�
��'��R�s1�#S!��TDqZg2�P�f�:t��L&��}��id�1�R0j������㣨�����9�?NM�+g7ѧ �rTln�+KBGˇ��g�?��־u���g�J!rS
�P��6�N| �8�4���	�<̻uT-7�,�=Ky�r��1\�vc�MR�Atc�CU�|�h4�3�%��n����TQ�
�=+;;rݳ7J�><3vИh����^�"
k�g ��ߘS�˻HL�����ˠ�DNjG~V�5�$�Ӄ��$=~O�� #Դ���|k'�~rI��H�� @58�'���H�7��D5X��.L��<#��1�{u��O�$;EoY�����v�p ='��D�ͅ��K �: ,�̟6�Q�����kU�xQ[Ib����y��L�2�Jp�6t�EM�,ޤG ��D*��Xг ���\2����U�0_x�>�k!�k��^�٦�+1�t@�����:PH����S�
��L�Xȗ
9�Iv��n/��0���9y�ΨW�~igj���ƌ���ޮN����.vb��v�SE����?S�l��.�(2/��?m��B���e|������+�ԫe�0�A�{SNo�Z�l@��Y"Z����^�4+/��9vE�d������F�R��a�i�TmmB
�a���	��jt�dl��Y`$�0Z��e��7r���7���JP���W���&���>�X������aPPEv�2$��-61���$(�k���D�.�ӼE�9U�B/����=l�Dv�0���p6yk]��^+�-��x�P��$�X=��}�YS���a[7��`�5x�>���z�s��.W��]���b��;I�G$���/��RU�ئ��I;������+��?b[`��͵�|`h ���={�)��#0��"��苝+��*�7�=�'��;,�
$@��b���SC%��$�y���a���/Mփ�ц�d�e�1 賧�	?�{O�zh�O-:BU���Avı�n���GW�5ێ�XO-����/�M�A+����?W�ޝ�OU"����H� �o��ؗ���}Ҿf�}8@�ӅP=�[QU+��������o�)�pN��dEka�8�64Ih�S8_�.�Ҙ��HmrWtO$#;���MQ� �;�1LL�����OFys��kZh����L3�Ľ���}���K�.�uX�#� ���^ޣv�뫎4v�����Y\�����G���xC�4����I��h���Zwa(�.�
:�6(.:p�l��֒�ry��ϩ0A$�,?�۸��|%?��[J�<�M�i��D:yvJ$n���>!� ff�V��X�7��֝�"���H�NwI߭Nu�/�Q���:�A��ƀ7m"�n��J<�3ވ��ڟcͰ:��?�c��;��Y�d;����Z:4�v4�Ny]��]. Au���0���yg��-9G1�6ej��!�s/�p'���Vp-�������y���?Cj�!���%8ә�W25����[��I%P�ܾw�&�
j>?��8S!~W��n$O���j�]���nz��d����p.uQ�(zɁg��>���O��Gg�TWH��yGl��L��̞IS�B����6�>�����*4�;��> �^�g���}g��"D����| ށBz(�R��g�*��_�EqU@�㇕(����f�9�`��<a����oPb������[)NG|־"���*��+��-F��mjh�
���@9)n����g����9����[ԭe���۩K֪�dV�����o{(Ic��I*��e�i����@kbC�o� �E�|�>���&�2W^_ҡ��:�����|��L�xFҬ��	�<���}�(��H����eO�����]�c=��Lv.:ClA��e0�F������"/�=a:�C�c����L�S�o*Ƭ�~k�K�lU��/��!�8�q;�j��s�o�f%u���B��%���"wj�,�`�I�?�mg�%o���1� ���xJ���n�/�ĴA�x�[���C�N|��^�wl}q2���}xxO\���ok���)��r.���}3ө��HK9e+���4�JH�L��e���>��Y\�cV�Rpƚ�eV���d���<V�ĭ�3)�]L
�E����x���<5�M���0��W�ۚ��MA��li�1���6=�+�<�gqF���#,-*ti����l&zӛND������s_ʈSnb��~W� ��$|�"<9�OP���+#^��X7��\�Ή5�+p0ڂ���?�Ec�Y�����0 �FN��2�bݦ\e��ve����i��6ܵ�+(�&����EV ��o5O�i{˥+Ne4���@Љg٭��/v����fɴ>��F@v�e|e�v�sv��6��++�#?h]�'�o��V�)%|7��r�X�#�.+!��U<�#�����f���������A)3�����<n�w���~��I����}u���e�u+@�Z�9~+���B~� ���=mM������\�=w�a�.S"5_!����Vu�y� ��Q��Wݓy+AVT�~%S��"�:=��Eb�9���Q.�%F�.��aKR��qͶ�z���������^��졞)I.+4aӨD 	��'t>5�ᴕ ��Q���rGb�����T�e�� �4tD�,���~��a��8��U�����!D�r�;�Ts�[.�^t�X�v���G�P,.>P-�[�l�B|�P6�N�r����x����$q,��O��D$�$��M����C�s�����t����Yʤaz8bo2����X���7��㌘$�M��R]b��v��x�ZA"[!��G�� b�TF9O����b��+��@n�nQ�CT��\�X�b��0��p����A�!M�Mps&�zz����	o�/��e����<)�z����+��t��/x�ʮh�{�ˌ��0 �X,�U�o� ͠`1b[ϛ���+r�?~I�Tnm.���qǙڂH�E&>�=��K?����,yq���~1
rn*��Z����&{<�(��A���j����`�zj�CO�XlxVHYEB    3981     4d0x�r/�P?^1o�d���Z��\"n�fſ���L�|��u2	ϻ���9��u�y�j~V':+�$o��1�%�Z"$ cp�?�9eJQXC\tw�4���P6��!�dT�a� ~S.�C��� �C�0�x��gY�0�/
���e�r�ߠ��o��O����ۜ��Y^�0��-���P�4τ������Hd��)O��!F��+K=�	��J���"�Dҙ:�����b!���u&p��94/h3I��cl�� ���F`���R�J0[�YnD�o��Y�,�P�Z�DJ��;b��Fyml������NI���"���ӁF��z˟ث�ݫlؚ�� �'�j��"�K�=7	�9�%� �Z�L�P���=\���Hjw� �j4�}��ۋZL�I?�݀�ʩU���������=������[3oN2Ģ{q�Kj�k��<]�tdR�}�	e0��q�nU��/���Q�bw��j����/���	1�@e��� tIϴ��.r��5Y������'*�;�q�����S��~�*�3�Eԫ��-,���
�L�Wkk#$峘N���Ro�T��ី*����c�$�U.�
*1s\�HQD��{j7ɭ�����1�S �9u��wbq�>�v�]�2�����2|I��D�t�;'�6��	 �j�&x�uzV����H93�A(dbǫ��qL��p�dD��z�M�0=��PvޏI1��i���z�T2����Q���&����+&��J�iH�i�&z�+P_Yco�r\�Z>�W��@+ZC�����Ǽ�$RR7��C�N_¢����tj��l�Y�NR�D��$��K�P���X�{�G����2�n��1��Kt}�Ɂ%������'�3`>�\���8G�x�{�$�i�����P�f'w�yq��e� ��b�3�z�-{U�����	8���U;�s���Y��?�������A�?�������_�G~�#Y�����e��N5������b�x��\��d�)t;НΗ�17�?��a��z�~Ico �X��f�-p=GbqQ��t��LƲV�(��0��^l�ս��A����õ ���k������r���CWݿz'5�o��L�↯�4���dWz���gtPN��a�h�v�k`��ፋ��Q0+��L ��2>dtͱ줥