XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��-�x�މ��QBͰ�h ����g���o�g�	ua�ZX�pDF�S��fA���-��H�zC���(B�{,+N�@q6�F�g�%d7Z����Q�{9�䌏H �z�ͦ+��4�~�$���׊C�;�9#THr���*EuN���[�v>��T�Դ�^�e����NC�S��Q�:%�A��J���V+�IjF��IcR(�~�B�� X���Us�����Q9G���~G��v������0�	|�Y�e��,��%L����`��L�ԅ��p	h��������w![��&��K�� � %���nE؆�D��Yv���������h��/�v�����}��[�E�֧��9�މk����j� 
� �w/B�O߀��<����������f� ��Y�@x��
�>>�\�3��@!�V�95� ��3n��&��ˉI�Cٝ����%���6�L�j|�Af^2a�io��&��Y���b�֣V�i�cp��WK��*�ö1F���'���֓'�1��̶A@1���{7��O��r��[D���y�j̇l``������sG��aVl�+����=���F�ѝ�&����}h��Y�������_K}g��9U:f���x~R*C7�T�D����oM��Uhl��c%#2��3�cE�]�~��_6�J�%���m���7Ph0��k3ڒ.���g�"}=�
`w	{�'N�f�{�_w��|��θ���u|r4��f��ĔnI���������
�XlxVHYEB    2bb9     ad0�'C�
(�W�7��������ܴ�H������z�z}�<͞�� ,�l�N��mڿ���L�=��p}#hƵ#秼~O���ٺ���i �'��罜�MN����%��sKY	�C���L�F���Ͷ $"H�ʴ�^F_�vss��	
ܵ�0'&.���签����|J�ܭc��T� @a��Wi�'"{�PE�?�z$&����^��A����Fcy{l�uM���lESI0(2�=��w�6�-m�Wv/�H�H(�p�8Z0����eH�H��w3��3,<���8Ea���K*����+ �~��R!xa���ť�$T-�}&�}m��YG]3��2�:n�G��M�[4��t�Z|�'{D��SH��ʹ���Q>�Fn���Y��]����yh��P�����(&>;�YC5'X�=r ��t?�tH�ˠ<��w��N��6�q�����ɘL�~%�{�0~�0W6EǇI��$H�T~wQ\��۴�w�w�>�%����H��_�ޖkɷ�{F����⎫�9.��Ly�C�."�.
z��O壬��^���l�:e���I�2C������U�tVR����C�ʏ�8���@M���>ۢ��
&�>��W��L}�����Z��:D��?aY��������l,��/�[g��#z���]�--Lc>NJ�3�(��͠��o�TDԹ+�����a|����8[o�^1U��臮�7'8���PL��u�5�o��N�8;����y����z;���B{��.b^K툇��~ir�E�a���(9 �G�NH��W-�d�Ĥ%�(^%�l��u'٬�T�	�o�3��@�8��/C��"�?N�"�L��fUS��F���]����9�(�D3fC��Kr�kw-�d�����Nr���2�*q�ߺ�9�|��[r!�g<��Z+��`79N6�?�We��F�5b�PaIF�͠���հx�4ۘ;έ%�aJ�M�eʚ3��^P��}+����<W&�	�����y�B�γ&���tB"�,U)Ϧj�����:��������u�]��@de�{i)⮄m�ơ}�"�F3���=6���"i�5N�)�z�J��5Fdo���}U�=���nꔎwY�j0���	v�`pf`x�����
)��qY�V"-j���|�� �)�Z�!� �����@D3��p(�~P�P��C�7D�&��-ƷA��fz�����6�۪j��I���w� U9v��ff0d�q��k�8K8��d*��d�Ώn{o�<^����1�^'�ͫ�]�'�a�uO��i8攗��c$(#��Lҋh:��#qՀ�h�s̷Z�t,�͇#�	��-��k�&DLx���{f�B=���!׾/kF��ÎQj�{����2A?�Wx ^\�[�#��,��C��Q	�#�%>D�6V�wF;)�Gt�ho��ªg4.�`QS���-�k0R'�:r4�1+�y���G��4�~̗$s�5,��Kv~N1*mԝ�$�=tkg:*嬥��;��?_\eI��qo�������!m��&��@s��M:¸s � m99�>�o�A�Ѕ�^����8{3�X�L=|����iG@��֭#������j�E��ֈBA���m�.�������"��xG���r�D|!BU�����1����*g

��k-��.��4�J��T�y ����L�"rB2Hzq��=Ш�k<�V����w��.�����;��l� V����(D�,47V�#���qσ��u�U���&jn�7���b���H����Ƨ&���N�㈉�=���?i�<KZ����G�7�Pj�j_D�%�B��08O��7P~M�M܅�`"*Ʃwg��WNN�1k���v��rh�SoK�o��P�����o;���,����EE��RX�m��>����kT�0��D�uv�~��G`.���)���4�0%�&0Kg�isr �_Y9��	nV)|P<8�!��x�DxK��;�tpJC���ct-��f�Ld٢<ly��	���u��/"�[;�2�+���<L����Zb�z�X�9B��!��c����íu�I�ߴ°F�,�a��	ﻧ�l�mg:J����7�?�/� Ѓ��CgE1}���b�" 7L�>��|�2|Fe�V�x�ɭ�m�@Z�$���ˉCڅk�зd6!��D�*8�.W$Fnr�<Hmvd��I>�o�)|� �淟� L{�3Q��hN����8�H��S5G3�	�\_�}�#m>#v{H��S�6-	W`<=,0�,zcH���G�3R'�_�"$At}ڤ�uQ@-��2P���O��➠Q�I9�߅e��2���T��N�k���yZ$ޣ�W�Gfb#��qt+Vw�h�����5Xd�p�^f1 �t��B|\/<b9��
��EV���λ\ܘ��?���O�����N�w�7��*'#�e�P�W<�Rxz%�U��<�=�x�]���'o��ܣ��m���48Sǁ1����֜�3�|)/7kV�6 �
�& A�'�q*C�c�A�w��DƷ��PD@w^�|�,>���C >Vzm��t#���@*��4�g@Vb�"�+���~��i�V4}���{���#tC�2�:�����)��
��q�K�:6��K��$����b@m�3EhR�y���'n���ˀ|@q#<���\��h��ĵ����9�+I�vK�8���$�xi���!kucSQ�Lo+=