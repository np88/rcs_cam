XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���p��,���i��|H�_�W^��я���(y�3Q��?��!��w!���q�鶈�{�����i奛�ku�6?��.���xR�q��5[r�T022m�t�Z�e����iϞ!�����-L���1.�zb�wmjs�^]A3�)�H� �C�jm�x���D�^�����0����ʸ7C��j�@ic��_�SV`<ƣ������yڥcꌫ��*̩Nk��TR�[�����kp�6&�n��_2�?�v����ꢚ�����,�É�!4/��Id%���ke���!"�e87�	�#��ɑ�b���#�\���W�3:��|7�!����
wB5�#��YV$�l�E����;��w�\��E7U1V/�k�.���K�լ��op�;��)�e'ׯ.KU;����sdZX��$�M�^b
���ߪ�hLciLj���\��X�n�e;+���Auv*'$�/���w��	VXۆ^�s�^��v�>���d_>�捽J�z��E��Ω;4���da���?�ʠA�_��'����b_�=\R/im�Nhl@E�P�!�MuoK�5Qb� �t!�)����ں� <�؇RUW#����[�n�5͜7d �%Z4�#�2	�^(�cAp��V�,f�X�W��	V�]'�:̈́^*�!�%EIG���#b
�π�]�	��=`�e�	������o6<紼�~��y�B|��9�h��^^;:�6t�Tذ.`Id��z��3i��i<���o*y(�	��XlxVHYEB    2df6     af0zhvǺ�mSP�ʤ���<�����+��t`�$'.�n�8�D���p�V�1�8�T�}�����D����c�����QZ����B��2�c7��)�tUdί5.�{8+����8:5�?K�B�
,�~h ��BVy
��9�_�2��8����^���a�=��H6�&'� �q�^�j�igeW���q��|����v��;���JH���QdT��� W43���E|T�%g	?}nVEh�?I� <z�"Y���M�e{�������u�I���#��u{A�Zx�u�g3^�]!"���;�������C5w?�MB���f�(Gcz��sP����4��1���� t�X/(V�>K��ؓ�v���u�Z{�t��*���#3��f>o8^�:S���V.�3|v�m�'�
2��GG��e�m�z��:�و%��"�ruS�]����Y��R8����F��!�[�I"f��D�6Z���i �8��rf���({X�&���*i�
Д������{7�n1	����ڀ�(?�����J]%f��p;�����aϞ�Z�m�fN��ǫ�n�|��,���ָ�2��ᾞ���qmU�dJ�|�\]��� �s���D�NC.R�o����e
/W��1���Zw]<��s�=X�z��#r`hGڥ3����B��a.�ԈTf������"�k��]9v���~�/�+�KL:����9Jي�V�u�PEbn�3�建�j����̆D[ՙg��v�����p�� �A1���׋�<�
�' ��Km�6���'ȋ�H#�oq\aa)����_kp�7-wY$-����&�R���7�R�$�Q��u��r�t%�^�R�\�A���º�DE?����u��*�Ӵ&��>W����.�F�x�̱�|3��5xr�==Z�m�Nr`gGC�_ԁH����h��͋a��.)��S���I|��a�(fv`�ҏ��M�������<Q3;(��]+i���)���$�e���05]�\�ɒS\7�����3	c.1`_풟]V�D�x��x:�+��Q�+�uL���%� o+ �<���{f���o�H���_�=�T�^wu�H�Bz�Qrr@ E�����ml�.`;�)���I�t��l�q�����2(�{�~�L��û�)��w���w�}u�x�+����(�����a���p������7_��;�I^��1<�i�DN���@�1j�:.Eo�3R���O|O������[��'�oS ��v�)MFEA�]���'�G��	=�"j)wv����^�Oq��;i+����Y�a V�Ldk��ڑ��3�����%����������)�I�! �&>�t�X�������_6`��q��7s5����u��0������eh�}{㫪M=�GPo]h�VH
���n9��9n?��e�D�qz�O�m�J�R���n�o��z��W;���\�u���vH�?���q�g�~n��d�#�ҏ��D��������5�IG��s������ב6q�jbƠ�OjUb����jf7�C-���Aچ�/yO\ <uK�|P��h�� (���Q�`�L��A�6ԋs/��i͗B2֠|�lx��q�g�O��y\�4���g��w_g���nJ��,��I�.�3���b
z�ѵ�M�n�hK��52&ni�瞅�>�3�ϡ���+�0��`�����m�J�/�:]4�w������	�Z�TAk+#��x��{�j?�O&���1*AF�[pf0H_m�ǚ�+���38���7J7_��L8��=[�[� _c�������V�>�U{�Kc�l�v��Nh��Zz����_�m��#S	�9XN���Q95V�����Y[)BC�1��A�Un���ȴ�g"~�U'0{L\l,��p��,��%C%�s�����tl`&�����O3H��KD�i{h�uz?��mhk�T�.2�������٨1��*ޮUƫm�z�B}EG���ֈaL�[-�M�;��]����Y�GP�Ҥ���ȡ����
o�p^e�þ�3��>Գb�g��y�T���<���V��)h���Ki	`5SJ.��EQ��k�D�����K��딲!�y��*g�8FLwI�mG\��s��y�rH�u�L�i�xzS9v���@����V�Y���!(���B8A�����J�P1"4�G�6-4ǧ���n
Ҟ[�� Y8W{�j�y��?��B�.ݐ���SC��$hsd�):��$��X�d���wB12��E��e��,�l��a�]��	^;��f�q�I��6y�:Yo|�G��}��ջG�s�Z��VjWzDV=��n�m�� @���'@�tպu�Qi�k�bl���:y�8�������I吉B
O�*�ǌkݰ�SN{�Ǚ����D��ꜩn{���B�d�=Ϣ�b�l��l }��;��՞E�ح�P����ݎ�o1���}����	����fX��<*
�I�aS����գ}�n[3kڮ�m�[>���.�t;n ���HEǤ#��4������ ��֫��$�'�I�7?�֯���@Y�UMAT��nۭ����w��&N5�~ι �(B5��ƻ�'։�а`o��ϻ,o(����2�8�N3�z.zJ�D=��x	��H�/.��������Ǹ2��=ʚ3A�d��3 ~���R�����R �L/T�n�v{�5��16_�G��n����J�C�V����P