XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��1j����ɝo�8~Γ�9�u����������|���9�T'��'j��ֱ(	�����U������Z ����#�^��%�d����I\�`����>W\&<�B��Wq@he�Z��É1/���=�;� " n��|�e
�-�"v`(z]U��ｰ��VMd1���T>r u�����w���!;++�H�.�]vOCۉ�����g�>��ŏ�bϦ�;��=�-e��nMw$a��,��Ex2�0(���v9��j}�DՖ��J�3Jq��	�t��̛��r+��_����7��A%]���I��Ѝ+L�B�w�P��j��Z�
q폝+$?~����,"��'��o��.12�����Bλ�gVЂ5��Z��v!X��Ǎ8���8���<ٕm�؟ˢD�S|q��'��$��V��i_G��+XI�GR6+�����x�v�t��Д����=��v4�j�JH� qVD�ױk�����k���y�=Y���U�Dk�>�c�]����6m;�I�ؔ���!u����[�MO7Q����<��o��^"Y��F]�|՚���<y��aQl���gp�]ٴn,�`h{8ӵ��:^�Ͱ�G��!�n���<���Ƅ��Ħ�
��Ӓv�`ş���dY��r�l����O�ew��e9���+�\�k# a�����P�������$J.K�e�h��9�D4�#��[p�s�W��F�;��#�ެ�.^j�R�]�γŉXlxVHYEB    5389    11b0>�k~�ѽ&����F;9&x"�x�����Gr=��H�f��������a������n�+�H��s�lL����:�I��1?S�� �h붌���l�ݎ3<N�,�A|"7��Eov̍�4��E�o�zP��	5=,�=^=+q2��4��2�*������~~��I�����Q>�ˎ�㏥�xt��L������XP��������f�*dxr_�՝���}�����{!� ��<'���<<W�/D���Ҿ+ṕ��
�Ja���A8��B���J'|�4D�����N���A:�(�����ڎD�=���`��p��Y;�Fp��-�����\�JQu�!|;��i�A�����7A}�R1)h3��_�\�]�0�Sg�Q�Y�uL#�t'd���B� ��:R���\�>�2������+k�o˚������?�{&�}X���$z�!���W� %�L3M���v�&D�Q�]�%b/�X�H6O�K�7�?������Ԑ�X"Ls��)ĸN�}�Їh�:z����[�8s3�)UT)��Ҫ������
�9��z?�KCaIY��w��ђU(+��n��[]sI��7K�i�9f<�
��s��⫙4����z$r
E(��3��t�3je��8��������I%Mx��k�t�_?��x\��8{0�fq[3�%�P@�'���������ݭ�����/r�;zQ1�`�M����H�C�����b6�ǻ��ϕHQ	���L��H,l��&S���Ҏ�F���K݌�l����oț 5@�y�׵���Z�p먀�͹�g<�?J�=�{>���p����fm*��C��P��˳O��+���"1�i�"��|��ҋ�vº^>���I��
�3����#��A �q��M!߿�#a���E�R0��E��=6F�yn�U�3�����G���`�(yP����
�5\��K�dx�
�q�a�Q���M|1l���$5J�	o��g}_D��)8�`p$ �+~+q�ȭu�����͉�UG0@�M�)���Q7�rf~(�[�X�LuMv�kHĝ_%�iX�9�'2���Q�w&(����X�F+R, ��õ�H ��Ǜ�m��S"��S*�A�xJqڲ�UZ@e
��y���(/E.�/ii�~߮����P3?S�Ǵuj��'�@�@�{ʥi�^�Ae��šZ�&,�R�C�a�
�٦%�ja�]�T��w<��}�;qc��x@y�MZ�;�o��ʓ��8��@���lKMA�.
2�@�׳d?�3�a}��F`5_N�3%�}�.Ϲk�G��+�S�t�]��� 2�@��DMtcF4,8�I����m͋����D����E�=����s�":��=�nc��bM*��}�>p@�:ڽ�,4�0�͂�⽍<���	1t\�\��&b��/���J��1�i�UQ�	ئ�-)�1�M���!S���,��'�I5�ʀ�w�S#���I@AE�Q�,b�10w�?�,�?44�p��NV�~��:4.��z��kW���{�i��>�t�:Q���J[�#�`��%7�\1lN��w�,8Ϛ�4\L�E ����싣�Wl��r��c�� *�ϣ���9�m����3�7�Y�8Ο�3v�}S]E�2�������~�*�x7F,u���ooMdG�Kd2`[������}ק�#��8�ߚI���=�'0R��:���o&��p �Z���(�͜8P�"<���2`$�F��Twjw��{�9%�=��������0q�6Z����-��z�+>�"/QN��b��EW����A��WՋ1ϥ{�!9�m��\�a��qn	W'�i���7��(m�̈֎��2+���EC��!�M��$�(Y{�s��t&��	���FY����`�	���E�N�"y�h�$#���cAW\�[�����2��v����"�w\y����Sgj�H1��%����%rR"�QSdÑ�?\ؖ�����j���xm�|@<���O��2x��E����2v�*��w�$]"
�d��Z\��}�C����7��)1�w*�.C9n$^	w��Ӓ����׎�A+�O�]�u��d�F��	��賝���L��5|��V����?��i��aV@uC�Dip�y��ϯw���Q_� ���O���&�y|d� ���^w̲��\���h���1 o}��2���Kәpk��/����>(�Rf�L��A|������c�E*H�G�*X�*����aߑ�|7ӀZ^��'7�xV�)����h?�wU�5��t6��I檐��{?6w� ,��m`��X�=��}� S�<v1\/�@k��?�=������9sZc��w�2�>�#�j0礖C�#Xg��2���"ݚ|Q��ӿ F�3���i��Rv< �fws����C�[Y�����k��.���yO5��k;#[�������r��h��}�']�r�F��L���4UУ "����43�}�q�(�B�ݪ��3�]��ε.��5Ғ���x��K*�
/�����|a���r8�+ �.�h���䰷�H�I�������@1����oM]t%Z�Q�� ��'T&��Y�]C�^�P���'PEI�LL鍪��H�ɢ�ګ�+T����a1�����Vf��f#8�
��7h��r��[��&.��y�@?�=��2�[~� ����'/�������:�	�]\���d�0E��j�<oB�2���s�D�H�A�]k,��0F����)Պ�]���d�M�B�qUJ1����c�� 4�j
�4�v��.豔mH�?N�C���}�Y{XNP(��r���H�q��0t ?.�#�(y���.=�j��pz��K�jPY�އ�g7p]X�7�1w����A�B�7��5�]h��o1Tp�;�UT^�ZpZ��� {����=p"3�S�H!C7�(���>�m��:���2{Qx�'���V�!�Fw�N]�.�m�Lh�UPk��Ǒ��ZG����ł��*�c��/;?�>���Q�4��T����.�2Ə�):X�x��	Ճ�Q�Բ�jx7$bϮ+�eL�v�vl��s��n�g�����d���B�-ü�s�%;n�f���;�=u\9��L8�ixX�iN^�EA$�iDn�&��N)�[kq� &	�e����l&6�� ɼ�>�����>��]��f�����Z��,��͜1ߛ��&1q����tK�x�nÐ�̇�r-b?!g��0U�Ll�iI+���NmӇ��"��kͣ��}?6�]&�H�mI¤Y!;�?*����93�,H��\�ɕ��UL��D-���q��(n���!$����+���E�B��H�g�j]�<��J��Bk��2����dv�D�K��F끠<���ؚ����w�A�G2�?�S�PV[��`e�G\[���ZS���,=��~L�!�38�9������}�D��m�\�f_�Õ���f�	IP-9e�4��S��t}��*�5�,�QB@�7릾��:Q%!�s��=�T��6��Z�=D�]�/3��#��ޱ�1Y%�A�\W�_��H��|xe�����.��"���#��Rh�&� �c�5��i?�n����Y�Ʒ�>�k���
���DC��c������C.!�����"�|9#�_�i 唰����Μ�6�u��������	A� �2W;�N�r���'�e����d����[���ċ@��(�t�K��=Hp�"U�#6E%]R�@֕�2a��V�l�geW��ԇc8}n��A����?ύ("��݄�֒`:��8�\ ��Z�.�-Z.�uKfr��>�el�"�E�'[m&|D��[��oS�9?'$���Q�m����c���PZ�88z݋����3��۽r��2�+�@���[n�.�\q�^b�� Wu@΀��Ty��uկ��b1:�w �)�Z{aM�.GV���M�=kc}Y�)x�dyQۧ V*��ğ��vVD�r|N!-��jMS��2գT���C�O�?���/=#>����t��Ë�
7e~�o:o���ʂ��M|�8�j�3.�1صSO0�Kɪ���H;�ƫ	E���M��(\(�%[�y������˧�~̛�U�bvM���#tl�Pm�q?�f �tt/���.
��+}+B����E�4��I�1e)u�v��~^�WzB�Jno:�/����4�����Zi�W��^�I�q��Ԑ6���#�|�WY��������0�叫�^]Z�a��@DE5}�=b�}%2��39ʎٜ�ŠO�>�q8�����1�MTa��W�rZ�@(k�V�
�n��{��2[0~!����B!jy���}��phq8��ec��=�F�'�rYH�W�!y�˷bg��"g'٨L�?�Qcp
��%(�L��Ϧe��D=�K��iy6