XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��vdM'�C)҉�iP�s�O��╤�'a=+�#�!5�ڲ@�@�=�o�����u4�n=�2`�3N4{-�W_����Q��l �n^ϥ\X0�5I�H��>j��'ȃI�M@��'������v���	ƥܖLIy�2V/q ;�n�4�e�5,��}����[Qr�z(��[�hUPk&-:Ǩ��UN�M8����m^A���N� _}��2sE���|6���"�&��7͟�n2��5꿖�3Ǡ\�K���5ȧ\��\�q����;����Tdd���b�7�á{KvF*!��~PX����
�W�.y���޻��+��O*�׎�a@.�U��H��n��wZ P�9�r�Cܨ�*���%�/�Ui�!�T��!�̀O��ӆ���*�ҵ�>z�h��O���7-��,ѴG�6l���Ez+Q�S!ly-g?�{������~ǲVL�� P�=��w��r����� (�]�\�-m��K�Q����+ՐXIB�����ԏ�*0R�_���D�\y�("d�`S&�m얕A�=S�	���n,��N�#�p�h'߷<]e��IQ����g�R�6Ǧ��ߒ��Y[����r�����{��b�ԑ���0ĝ`Dԯ��9�rn�n:?�Ć����3т7��U�aE����M�ctP&I\"�1*�����䅊/��Y6�~R��|�u��1;s�n)���#���L"r��A;��UlY��ٍ��@�(n��
O��8�տʦk����x�[d�T+;�XlxVHYEB    3d61     ed0�#�Kp�kxf<�Iq{�kk��Sˤ"��_��,E4�4�ӏ�P���\ѩ���Q P�F�I%怴5�$�7�ڊ��0��|�dG�u{�gE�7K�x�'�mѶ;mY��>�U���6���4S�^�c@_b�]_�;���ʶ��zjOl���ܵ{.�L�$;E��������`�����6���_ѓ�ReA�~^��:piy���2G�2|G�f�y�+�y��_g�=y��ps�j{��b����b��#��Z�t�� 6�Z����|�"�����D��l��	bJ�s���>�K�y��Q����O��J$"�ӕ�qp*���s�2����S>�����l��i�� >�b_��ωoo����W�^��S��%R�Y�''���V�:*c'�1�\���7�G����/�&	��[rD��3��o�4�|3?*�S�ʼ\%� �ӹ9�%�Zs�+�o]"�G0�u0�ͭ�p@�%Z�œx�#X�3����6l�z�5�KZ��N�)qs��8�i%Ľ�a�����H������r���m*^3�Gb��H�Yg*BǶ1k5�t�֤=l)A.��c庰�F��*۲�|�U���Y Y����]�)j��{�z!lM��%KM1�2=W���~Q��ܨ�ܬAo��y��7�\1�'lT� ������#�����)�����:G�����a��p����ͭ�)eq�Lp�n�K�P��:�R©wd��и��8\������np�'
�G{`�;j�}�׆IH�C�$Ki��(�N b_\΋�mKTJ'��֙4h��Yt�;�{Ճת�8��߀��Tp��<���[�x}"aB '�!ԏb��f�m��+�Ԥ�r7Ig�Z���X��{����
��`��P�N�zf���Dz�D�^�7�e$�P6t��G<ɲm� ��r
��+ ����q���[�]��yx�"n?��'�h�o[f?t4Jm+Ly\*�Ϫ4办���e+��EV�
PvU�|C;���ϝ���$�[c����F�^�/al��+��$�Wq�h6�P��oa�-����� �^��A�*a�|�)�}T��Ԋ�y�ND&pN$Vؙ6���~�.�4�8�W�� 6����Һ E��ql�M_�����]�쐧�u�l2d5!\�Ub%�P�T�p�2Tu�	6?2�먺��r�6��((���"i��alߡ�U�{���;��*&�������`[�u��W��p+�h�:¢���}�6�DI~��� Bvm<�Jٻ�jK.q��niF;������6�s1ؠ�(TX����L�=T
-��!åjY�����=F���텨px��C�*)蘹��Bє&�E7�1��FK3U���y|\� �hb5�^Jew�C�yO�L�.�<��p����E|���aţ��sڥI�EIr�ʶk��Bƪ҄�8馗�
�q���C�"��wL9�$�\�V@�k��8֐�ό�!h��9�98w�~*nÄa�{۠6ZS�%��'X<��s�K���9�S��T5,u�����|m�0Q�(mjQ�``p����Z����t�X���ӹé�l�Ԩ����J[}�5�XLǹ4�����7GW�ӝu�Fu&�{��N;���B�S5>���[�L[,�f,`��1��a_����'�E�yI�̈m���Ar�|TV��TzM�ފ5^_`�o��#�����6����Ѽ��T�q���r�<@w5�K��/�g�'����^�c>6���"K�'���X1i�`.�˝����*]fK�%?���Q��{�K{����74��A_���&R.��l���W�N� Ե��� GҡfO���F���lg�H�F!<�[	� �r�	��Eʦ8���1���Ws`[c��C�*h.��6ֲ�d(�4�k�P����e.q��>�3.��D=�w���Q�]�qF���J��AL��|}5PdRS��V/#-�0���l
v�:�O���&E:�B� �Ƀ�7Xꭨ᳜7d{%n����Z��d�w�g���+k����!h���Y=���f,%�ts闺W�#��d"�"_7"�?y�[F5y�h���P6�I������m�}��zd ȡ7�
a�c0��N�M3X���m��%�����g�HnM�86�T�<�Ȳ��L�NI�!�e��Id0���G_,5���-��O8f���(K��0Ig�G����mZ8�o�zg��V�v�� ����3��E$5�aW`�?�2V��m�M����(�P�\�=���M�]�ڙDL��9�F��O�Vrq�cpW��>C�����!k�(×Q0�c�D.���MLTգ��<W��B!A�O��C������Xx�L%��t��G}z/haϤH��	f��؎cڌk�k+7rY'̅��[%����������Ƞ*�J��8:�#hUP�d���ԯ!ZU��1�Q�J|�}�^m�\b�����y�t`�Lѵ��܈����8��A[K��ˎ��XP�&*Gj��.���p�j���F?�_4���_��jM�^��Kv�9��V:f����z�A�jt�_��n!Dl�-cٓ*VRj�3�JAxM7w�B�m�rlS'!��c,I 9T��Q��i�a��3=��)r"7�_���!S�2�zx��H�7�M	J �ψ�	0�.��*�5�cᮞ9�­���IfT�u�Pe|�3ɿY�&����i\��>�������?4hk�������,!)�P�zb��V���Ya��uD�6^n"=̎0�财!��)�J�#:�YT��߁��M�I�0��[�)�5��j�Ϡ�SE@!�FE�BS�y)��Ʈ�8.x�r!��"8�={$�x�������IA�*���b�0�:���*[γ�SY~��Ip(W�$ibi}�h�Rީօ�l�{ڶt{���.$����h������ 98�鼓Bbd�}�6f�p��[��.�:s~�_��4w#�!�W�=�-�� ����Ң�����
�.w���PIK/���X���j��
�QC���!��s��ӦP�-_�M���Qz�����;<Z�g?2>�����Е�J3U�Gp�	c孿��T�_<��)��&KGͻ����ݜ���F�#j�pb�9�k2b4q,g��Vɚ��D�.��oT��GnQ"�fvCܸ}>c��.�kU�`���\A��o�1��2!�g��c���]n���sXg�}���Ez^���d��|�*�d]BR�I�Ӹ�̚3j5��tM� &D��,�
M�,	q�uHj�-ln�Ց�df4��������m�4�_O�o�a� ;F�Ci���V��y-e7����4�~��z��:�H�ˈ�pޅ�:����wQہ��?j%�V+D!� g�4�?�,&Ҽ`�ʗ`����p'�|��5H���U����<��Ø���B��6��2Z������ �$)  x�dcT��R��O�E@�N#:e�1���m��U{&��i��Ø�IP#�;�~;��PW<!�΢^x}R�^��t���V}.^����-�H��!OI��U-�|��݇�%����AoJ�c{��H��0�'p�@tZ4*׊�ջ��F��=�e�Z�rcR�\�/Mr�9�����	�҉	�h�kdI�tM(����Ի����Rl9���'jN�������Fm�W�&>��Z�΍k�ha�44fZ�l�(0�0	=:äN�f7C����8�=?��0;