XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���$\�]���I6���2�D��t�2$�
��}��*�>�Z�0�Go�0pYBA�.
*��H|zkG@��HՄ4Qr}.zPr����|�`?�i���jt���kKN9����|�s���������j8��BKǉq!����v��g��/ј'kq|ȁ|���('�xmk;���D]H�S�}�6ƭD+[r���Ȯy���i�P-B_�Yf��vS���[l��K���QSW�K ����K����&s�+T��^��:�kYo�^>�ro��U?�K
�S��w� ����P4
�4I�����;v��������ԋ�@cz�u]��~gz'�{��X��b��Q|ڑ��Aխ-7i��A�"�O�tZ���No�l�b#ۋw�9�a}wy�R�ɸ�o�7�g�^�~�ܥ����}�Sb�q�A��������q2���A��"�:}��#U�z���Ia�q�� +�����?�@�m�%Im?�G�*�6���-:jPM����Ļ~��<������O�!�h,
\�W�����M���>7��Sjk�/�r�u��`v��%N��	� ���ߊ>j� 4`;�ͽ,�4�;�.[�'��X�)Y6���іkPm�{�X
�w	�������U��I���N?hK-��v �����*�zq!�J�nR77�XE{���WU<���*�sg�].M�o;�������p�654X�K4�����X��+��p,�k�XlxVHYEB    47d1     e90�,ԜJ�wLA��=Z�ݕ��#��k��L�O�摉��xv��QF�@p�Ì��=�9�?�T��x,\ؖ���Y`!�c�rW	�"=
G�H)�-q��"����$��È�Ys:���l���me�8��`���i+� ��skPy���5 �+e�
�3/"��H���fL��۲��a��t}uR!����-p�׊���/V�!��$��[�M2V� � ���󣵪�!d��kq��I�����&�vh0�/�ʏ��X���^�BA�_���gz�P�����XpL5v�om�s����z����@��/EOj����Fr��ؚV}�I4��@.�^U�o	�Z�J�Q��?&~��Ҿ~5�`F���CH���[�_�>�����;��I0�M���|�a�hx!���|�C��O��^��+Z0GG��&�UA>��e�W�]��F�;\&��ĥEO��j��M��(��E�z��e5��n���h-p(R��b]�'K�>�ν>������D�Bp���X��z�B$L��\�Gr�԰�b�b�[�,�aB�䰒_�3�ك2����a�f]�*�x��f��]q[X����s�'�bm��$d�ªb'G&j�'��3T7#J���;n�G�ϿM���������uP&=9�,��2�ِ���S��.f�@�t�D׬EO�q�w��ʸe�&|������ɫR� 8�����+m�e��<�l��DȗRqv�Sྙ�$#������@S���Q�X�GЌ�E�C�Ѹ}e��`J��W��p�w�B�f>�d��_�T�
��\�,��l�]��3��tߓ`�c�jIUDf�g�M&Ʈ�)��2��&0�����a�%#%{k�"�I��x�'v.6[�&ǎj��܅�Ύ�v&0�eTD(��!���)^'���S�����U�ㅫ:x�@��W�	n�Ӂ��e�7\��?��5��)ܧj�7q�-*�۱R{�-!�b�/\&�w#W9+��A�sTI,���d���V�n�%s� qM��;�*9�bL��А����,�{)�iC�ѳQ�x[���9������ς���A濕�la��~�&���O����h�e�uɆ�rg�c�y+0i4Pb2;���4n%CrM�9�{��D������C�/"L�3l�w����i��ܧ��ώ�ˀ6O���\Z��Τ�b8���{���M>1�'�C�Q�}�'�/��J/,���^@���'>t#VM�˷����q��L_�#ţ��;��
3{F����P�҆�8�;c�����ϲώ�`�\��%���{yh���x�ZrD��F����`?.�Z�$5�+�d#o;f��f���c	�����G `�sHb����x��{ ��(�r�&�/�K��KJ��c���^�V{,:��
��#�	�B�Iwq�-�)4M�V��ScG��Ěb�D�#e��.$��&)G,��
hr�S��VkT�<��mƗ���ǜjX370z���|�i�	�ѿn�p¤���X����/)7�i��%�g�O����/8�c2��%�4I7�����I�ښ�-{)\`�S�h�7��5w�����i�v�40$Kx�R�h\8�9[����ߋ̼���=��iV�_�j�$U �fVA��g�
��Wh����R�Ѣ���I�L�9�Q�2J��|��ԫ"&K����Eb3��6��P)���%�,�W�כ�8.ͬ�[�.�l͢r�	s�c\P!�<�\�V/�)G�Ē�HE�6�`�,�I8U_�e���C����^���S4�[�4��yˋCl<��bݖ�j��@�Y�����-��aB�^��S���$r��iy9ks|C�܀ɳ���˩�zg/��B�j(���qs��O��鯆6j��F�o���Ѐq�r��
���?<Ѣ0�躿o%�m].�=-�`3�r��P3�$��A�^�F�G{6�;a�T,�s;7�)��ӞyvOP��p���Dѡ����Z=�����F?e��١�&��1�t�F��ݓzf��l�aF'��,�
i?�;�t�) |�	�}�F$oE����Eڟ���� ɫ�[�����F;�ª�Ţ� ?仝�ވ�4���Q.�C��&�� ����;)��~��#������@��_�\�/�I}>$�y`�i�a�a��|[��9���	�����9�|r���f;CQ�o�J4�� o%�a�J}�D�D���.�+-�ȟ|�յ�N	w��$UVq|�VP����6R Je. �w�D�n�ؔ�;���8�c���Ѵ�@PpC	V&Iw��>R���Wd�{f�*�e�2{�	J�Zl��Ƈ��Og�k
��H�>(k$b	��~�u�g���M��c$�_��1�|i�>i)���_R?�6����]ĸ�BЀ��r���'����IZ�Ú߼м��]F����Y�<b��Ur�uͫ�+���(si|H/����跕�S!m
�L>�~��'�M4��8�~s��jK�܀$�Є-���������5��L��:�@�h'�'�����9�H�;������(�|7�0���aL�=��O�t�sۣ=�ϐ�|�dd���N��Z���T�n�`2klt��J3�*�BΩ����tDd��|�3�Z�>LV�����ڶai��&}��ށ���I9Z�чG�E�\&��ݣ�^z��X����×��<q�q(���M$�<V�fAY������[5+c�]dD���C���&������h�'7����j����7����
�(�� a�k.;���l�l$��x���j����w-�L�k�_Lr�n��~��'*�u�?Jk�J�WΥ @�Vg��h��zh�HvF�<j��T;�.�L[y� 8c���hT��d�����Ŷ�G`j�y�Xܔ�cPr�j?[�+�Fv��Pc�A��
���9�$�_U��8��2�o]�u��4��¾mt�ҞMC[+��ͬpjm���;�aY-��EJ��=X�J�=x�E��j�F*�Ud��#J;�[���3���s�u:<�� &;g�A�I��p6=Ό���C�����\@���t6�^�_&�X��%�l=\?���ǅ'��(��̔j����4�2������ߺ����R�[8���b���D��Iq�4[�m��DE�ԉ� �e���DJ�*�P����������X�s�ڤ����1�}�0��*|�T-�
XM��-�8
�Ep�+�Ǉu紀�(Z���S�Х���xNl�*�	������G�j\����O\M�~zWi&è��Д���o�<��VJ?O~������JW������vYQa|Kv�K���Wy�G�f���V:BC2��Q�yݽҒ�0v�%�����nO[�+�9k�c�s�\����2�
�ϗd���.�^M��fp<��!��)sj�P����$-Aw�P[����J��c�C���ïk�Q���`�r������N�^"U�K$�}��������?/��9n���v`|�(j���,�J=���� qu��KQ�JP�O�X��P���&�Bn�JB�B�A��wR��f�@N <^��]�id�>�aaI���W�����_jw��4�3V���>��7��=yo*�YX���Ε��0���2_P�