XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��"��6��Mri�>̹s�#D�J@�(WJ��,}4E�Oκb�QK�X��A����A��Ʊ	A^����<nT�LJҜ�ƑC�E�`c
	[Q@gsI��@�`h�_�9��?�^����پ�s��J�1[e\�ӕ>9��'�Vw���9�:Wn?�W��ϕ����|�տ��l����6/2*��E�!!z[�dW��)�����'x�ο/CY�@K�Q�W�+^q�Lh���-4���>�k���N�^<)�7�V��C�(*R��]N$čŝ�0ǦM��O�'�������fF��)"R���
"�� ����$Г�����8�Z�#�!�v3E Z5�Lΐ���Fw�hS����ab�$ƍ�!c+��~��n�'�����c[������E��hKƨ�v��,�.�[R��-�V|�Q�+���C�����g������L��y��c��e���F�6���ʦ����@Ǒ�jP8�g8A�*����i�d�[(K`kw�CX
5"�;�֝�J$(��_�}Qs��Ϸ�S��^���)��ts���B�Q�a�7|1�.�
�јMiK8��BP!��1+������{���ȟi,�Ac>6�
���a�9VsL��ރ���U^�2N�n]�����_�u����;��'.���iX�8�rڮ/��t�S>��\cL��54Fg�qu �Y���'�Y�ӧDf|�*{)pHV?�Fv�JP �㐈�-�N���Oɽ��a��0��A6�ϙ���;��:�' _�7��XlxVHYEB    c3e8    1d20���\�k9,K�ԅ-��lO��zė|v��3�WM�Hpm���8��V�~#���_ٙWH�����:�{N�nV��|��#�,��#�a�`>}8�qdK!���s{@�j�zwQ��0�b���y����b)��#VI/+N�:'�����=�������ȈK,����xj��p8X�����*z�n)��|YYW�W���S�6�;�<?$�~��
�N�lM�R�hH[<bB���2� �g�����f�����}�Ʒ��$��B(����AH��@]��z� �V1�ׁ�ŚN�\�qW�vŉ��'6��\�=h+�u��uH�b]������G�F:�N�TrL/5��ۡ��m�iYϤ��^B���e��e��6~�
�o��б��~Q:OՆ@��_/}�t�8OQ������Wq�£
���P��T���M�Ȧ�����"�W�6��^y��Kd&[}5���O��p϶^�٢����g���4�?r���$�N�|\�*����v3k�ϖ�Za�ca����L�5#�z�L>%�^�.�kTc?�m?�x`;q2C7��hn-�l���cc_1�('6���������>�=H�bR�ݕ�(�l�*�2ǶR���������@���z�c��ޫd+t$"e�� �$p��
��"]�	�Z�Z�q-��1�
�Y�	a��7?�8�(n�oVö[a��m�cS��X�ъ��4���K}v����� q��d�Sԩ�$n���S��fVU�#�=/�+���s��^�^/	� �zw��pi��z�%�I�K�|&AnC$f�L�+*�*�J��A�!��̔+����_� �QX�Zz q��D�}�V_�rd��E.W9��'�B��w��6�U��}��s��c���-�yy�I�Z������d~�}a�!�H��a�<F�{��u�*��(2V�ub`	��^.�}�w�~w��T�����Тd`�EΗ����%Py8���Yk��c�8��!��AׁI����imm9�Eǧp�ሹ���Ad*C1w7T=��C�0I��?���J ��;��������B���ј���j���j��0~��P�f{���0u˾��?���fu�"ݯ�J㦾�7���ډ�����PH׬����E&�tE5�{��3��SM3]RZ~Jp����B8D*�d�:��u�����K��>)~� A˓q]!�~��GTDj��@7�Ć�ѽt�|w�u�tCym\���ϳ7��%��b�J՗�����p� �ơ�LE�&p�<�ł��Yh��  �<�w�N�/2 ��MIw�+��1*��iF�����v9QS/�xs��7���`������B`����}�E7�sm��g�`��Ĩ�-�B�~��9�s�ӪZN~��\���cY��ؼ��bn
��-���s�^�Gzӿ�n_�E��G��c	*w�;h����L���/�M��y�y�i`��eݭ���p�+雐���$�%�]�*n�H��6z��ѐ�'�WM���W��8�XX2�\<��]�a�8�dO��mjj��n����6������0�����?���i)Q]���͈66k����,�E��T	��u__g�xd� Uq��YF���'�0��py�d����k@(W�#�
Öt�W�Yn$���2�aX���R�-�޷�1z�����ϓ.Kj�E,��|͊P�*���n��.������%��3s�ʕ3Ta��a85�^�rz�SPlm
2}�耷׳-Z9	g7�B%�oO�����7���$�noō�#[=��!�_��;�ӋˋI�"���y5��<a]�5��A<�e��*PG����M��QH(�N��<��� w8�H���7=�6tk�`0�4�zld�ϱ����1W�����1~.S��k|fÄ�˞�B�ȍ�C%���Rlc�"p*��z)�o`��u��e����: �E���m����?*w(u�pʧ=��O�s���>��ŠĠ�%���q�c�V���l�E�jſ9�n��߀�$�s��C�X��-֟s����ɸ��r�Y"�OԻ�0$M\�2�D2�əɶ�bt@��R��)�g�'p<�g.�%9i����{�*��@ EgM�&�C;�A9Jj֌�����5m�	�s7���2���tH���%�ؾa^�j��}�~nt�s�NMRKuX����	���G� /�����;��;kGӹv�����i0��,-��K;��\�g�s�i�s��:����]vW�옕h�YE��HAU�}dk�&�����l��UF1�����ڍ�Ӯ�� Ī��,�@��<�/>��lG��@�+�(#�%cX���l]�}Q�j�yz9�t�#�'Z�u����g��;?�
�LN)F�5�->af)O۰�,��D�6���6��^N��pǰ�f��i��x�F	��-�{Ӌz)q>D��W��<eb�o��6����x~�Z���ש�E�.�&��,��#fjz�&T�#9��G���~Pm�(Qѱ��94�\#׋��	����b�L%Y�70'�����|@g�����3@�A��E�L�y�UiJ&US������S�Z<�__��t���3bC;��&z8��{�Di�Z�i�e~��6�o~���hv_�JJ�ۇ`��{�d���ҭrIIw>i1VH���Sqң.�W�S5�tzYCU��ˊO�U��`�_'�� �!�*�T6��"F̳��d�F^\��Q��/k*hN�?oXt�A�K�0@Z%���ԏ��7�!�׈P�J�.�i��)�R8)�H|�LD�%R2��F��m��(��f�a΅~���<հ(}fx��R�ݘLe*�PC�*t�{�P��Zk� [eH��xdGO�h��)&���Y���u�k������ ;�a�j��z�ȵZ�z�����T|rs�BI��J����Ѳ�c���r����fQ2!N��r2�X�l(�f��:W�/]��O�dh;�C�?���7�I�a�j�5�z�e;�uܝ��2�o�P<�u�1U
��|+4�?+��o�㨄�5��<��3�&��^�$���O�>�y�*�#���P��$�4���Ք=�
��c���nbD�Ėt.��7��@��)Ph��M�s���q��̳AX�ʚr��bA���/Y˼��q� Ib�
�RՊ*mߣB���D6飌�@�y�@F[�����wX����ܼ^�֨er�E�m?��zzi��`Q��S���K�"3����nqi���>�>m<�'�W�/M�C�LP�:+������*3��������n��^.9��3w̮��<�"P�V:��}ZWo�جL�`�j�B�{���z/u�ˀ�FG��D7�óo��?��e|)��"�	����藙$��&,5�=�W�c_#��$��
�?�����1?X��W1����';
��	kd �o�DU��o�JH�LË$��A����<���e���h|3ݹ{��� ���ō�+�‒o��/f�'�3K���l��?��P���L�?��ت�Yr+;{�[)�0l�7���V�0N6�uW��v��`��!Gu�i��X.q�+�$�,�M�5����@�%��ZV���
˺�l�Q�kG�6�mc�I����@&H<*��7J�.����r<�"��.�p��<��P�l̇�0⺘'gs�u��_*¹p����rN�ϼ�;1K��B�
�R������5�	�[C XC���Zh���\HyC�a�Z��W�뙟�/�-`���?>�Y�^��zJ��M���o�S��5�%����cmu��0$��i��r7�#�b�>c�D�?r�|��k��8��4�s�)2�%x�n�+#b��\�¹Ѧ�.k	3��W7=z���=_�:��$h�@��˥�����pL��K5P�Ba!� ��$�b�=.vM�?�I�X�����*�ܤ�Ke7��q��TH�B���P�@�@.#��	>���CT��ň��n,/>�a��t����T%�6�x� ���6
9�����l,�Ҁz+ �j�����<�_p.�oH1m��E�h���:�SEXWQ0���a�'�%�W��@�C5Nə����I^!ȏ�؎�&Y��ĻAv8+m����������RG3Nh�j~z�Ul�#x��W����ALL�Uf~���_���Ű�#��5��wq�]>��a7'寂���=uwo�i����ݓԱ��	z�-�����D]1p"�3��#����	Ć����S}lw��U�uJ�*�U�{whQ�%s����q/�9 Ayw�x�H���[Y���Z��~�d�YKQ�@4o��ri���%O?D{H�P$��p��N���p}'�]o� ��N��O�#S�Ş���ƕ�au$z%4Z��Q�'��>e.�S�� �(B5��R�)C]jw�&�Tڙ�Y�[��9٦RXɴIF�����6E�f���o鈶�ם��
���^�Tϛm9c�ZlL����� ������%L�ƺ�|�Y[�I8�o���UU��p�{]`�p��H��Y���#��x���V��,�9������<-��B�A�����C��|V��:��婚�������!\�m<\�MfU�Z+��� ��{�z����M)9��j����b$b����Jo�|R���i?y����	�;����!�,�� ���k5�o*���5l��,�1��3#> ����
k�`�E���4�H�?���G�݄�2�ͽ��*�������Ҟ���!ȭ�1sc����)�oK��]�{ܚ���&r�A�CCC�@�S���Y�:R|-��*�N�2� �A]jT�GWu�A)󟦊ō�����>DDC�t�����Uc��G;�w�>t���D��$�U�݂bh�?]@�{5¬�+N��q����,S#k�t��&�X��l�v��a} Y�����ZD��b�LZX/����d�q�*f�XsJ�Bxm�W
Nꮹ�*˟Eu�B{.R',�S)u��$�3���zxp�t��+v��X���B�69���c�����ü��>�oo�G�{�0+�뫚%�	ײ��G��r�:40]��[el���?.�>
N��|��0mw�Wkw�8p��H�*=��rc� �kn/|'�+�¡x�^J�G"M�%H�+�W�� r�u���z1����=� ��åe&��q��<�c�6KW�	]�Yo�R B��d�,�[-��)�de*i��N	)��]�s�Y	@莴���.�,[��P� o���s�]���Z�J����l�2�s.�ƩP�JBD#FD�j�����%|-�O�`�0�s�Y�co���<҈J�"��h�'Z�	��w��.��S{��fp�z��ăLw��'R���%$��W;P��2�a���*��}���r��~�Q+|W�mOG���k��k�] ����Á���˟�z���>כ�'~��'��0����X����m��,�GUK�`gl�� %��z���"��!��A���t����H�$�\ۀ��W�7��ePX�q�z{�������1���gf}����6:��n5����u_tс����0_����_~�8��ǂs{��C~ >�r����қҎ\x�#\ �7��KR��|9J�6���O��~�2Pc�0�%�w�{�G��0f��N�A�qe��?���j�Ǽ
3�ě�U��(�7�o�'M �]���6�v�N�����pWl��G-����Yd+�z�cha��	u)���c˹�P����vƲf]��<*	��]�v)�ԩJTqn��r��Ϡ'�ꛆ�F�b�]Q�i��Y�(�"�p�$����$�K3��0�<�`�u��Q�Vg�h��� 󢢟'0H�w�d���f1ʲuXK�y|�W.����tN��ڠ��9be�Z��d��:�̲k�[��8Cx5ɞ$O�Q�h�r�'���"��vB�zYs��dVU��b��U��À��=
r��G� O��#e	=N��+�u�N}�Z/���ܚ�xM%�82�S�/	_��j��I�79"F�8á/�� �[$qN����	�m��W�B`�����%_ɘ�O,NAf��>�ȕ������(���S�b@�ƙ�?�:#AQ{'�Gy�h8�0D�9z�鑉����!��J�*��F^ �?��BE�E���c��&"b���Un�.7.3�D'[�9�?���c��=�V5|<g��(��DZ���*4���vnk	�q��H�j��7�٬��V��>�[�;��Ѷ��f�Gw�������E}�!�-��_"��N����A�X���t�)��r�:�E� ^uD�>�y�f��昇���p��r�9;!k{g/�ZH9{�H��(�)r��xAM��)�}Q!��i#�����G�o�5O9'�܀�%��+�K"i�L�]׿z4셍ޅ�L׹�bQ���Xu��<ż%w��K����M����,�(у_�FF�&��8�0,@	����8���+G9�ٵ���d���X�/�)��B��_���k��ܷ@q�����W"s7	����Q�߉���֍��8�|��	?6ޱ螯󌣜�V�}̨�lȝ?�����iu��`!{�Y���;,��L��ߓ�J�,�ϗ@��˲�3e�$I	z�S�8� 9�	�ɼJ��z�
����ה^�6d�&h��t4�b2Z-z,m�A�dĨ��H�)�G5�\�ήK�b��;�G��l<Tp_1�֣^oX���A�����/TY{���&�/Uژt?�""P�˭�������Oء?�O��$�D9	��>� |�f�d�X %]`4X:���rcO� ����io�tH��z�˗1����,��sRi��%x�î�k#��qMk�ׯ�.N3ה��CA«�ZP��.}d�8X�Y�M��#����t��1\��k]�I�6��Ϫ��Q�����xc�YI�����kq��T��P&*�l_����Ժ�A����ź��@����+}L�c���)>WM';#t�~ɸ����3+ g^e�~�����4�o���br�I����~HX��%��}��Z��H��(ޤ��gRIAF��b�\I~ph�sG�#/���?��1�vp�V���m�z��(���o!qn�����I���F����nЊ"w'��VL>*��W���>�����gVoܥ`�ۣ����m��K���A�l���&bX�Q�Eg��܎�0�S L�zpr�T�oĥ�9�����.�0��/֧L��
-fj�~��7������U��� �#ҋ�ӼƲG�y�e���*��u|-�6UT0|p�\}p���>"^�}���^���x�U��O���V��Z��-���ǺXq