XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����$��v�\����%�4_�3�<��؉5��W) 4)R �Y�b��f��_��	~�'��$���Ժ��6�ƒ�2�jZ��Q����A#�7&��A7�:�{��آĳ�i��s����우 ��ۢ��\ش��xr�\M�6�p��g��5e| np7!}����0 &#`�=70��'O�	�B���ۚe
�۞��]ħ�_�bL��P��-�-#�U��'�����ވ	p�"�@H�����g���z��qU����
���j�!�c�?<�5�o1���ژ���FyC����g��l(���>��H����S�Z��:��i+�8�:2�!-�m�^^~���s~)~rafyRa��@��E�XM�E�~�u;��dY�g3��\U�n�*S��]����݋���C���zcW}Dh{kM ���%��R��H�#^35�;q4;hE�].�0;=�Y�;�5��̧<C�x�O�FX6U;�������
J�4�Q*�Ϋ������p���n!?(�a�����mN\A����Y��P�.�����܁%���n&8p ֘4굓�1����T6o{��nK�������[�b�:;�W��'�
��V7�
Pj�,�~���|tZ�����C�Ñ�%D��3	�����rk��v8WŀOU���+�]�D��,פ�E���3U�T��g]�d GZ���p���h�>�]�&��H�/����-7ȏ{��
�6׶�p�w>�$A[qU�}x8��9-}bR�XlxVHYEB    1c45     950����k��d)P�*1��q��Ї��A$0I�2�I.���߬Byp\"���8͹Y����c�|@WֻR���c�mdR�L=�b%6#1�@��Ch[1�9P@4�J��ϗm�@�����U����H�.�ל��!��!������ 	��` ��X��
#���R�yc��7mn�g"���̺[�j4,?��m��)�n٘#�7��CL"Q�X�Fĝs�)�^�w��0�a]�ì_|2`h�. �1�t�m��W�E<�>�6}ւ�k�����._�:&Ɔ���;�w�u��0����E!���lY�p�`��("�4�c�)3�5�
h!�i?;&��=�W�G�@�s	�ѫ��\O[�S����.���s�� '��QSa�SR�gR�E�>AQ��e�ՋG�k6�*��f���.Y�����ֳv�kqz�vZ�UɝdO��6�D��T����H��n�,H�L<#`�H�׊�R�������2��?ĩ�G������PNu�5�͂߰N��x�T�ۗ����DWT׶��L�H��j�kGJ6 �_���\�Z5�J�}�a���L�Q�qP����n[Py��a.|��
(QK�������V0(�u�%$I�T��w��@�Q�C4�dT��D��:!y�ݲ��<5 XLt�k�7�GMZ�����B)�"��Fo�4���L[�����3�1(��t����������mr��(,j���� ���'Qd��Kf�*�K� � l�8�H��ޤI͐�3D���|D�A�(�Y��Y�F�;<w/�7���9^oK'C����긳�����.���+s�1�p�PJ�~�����]ꍾ5�WY����V� �{P������xxSo����o�d���M��{uyd�K��g6������E�K���d�=~H�t/�����P���\g�*A�Z6*��,��l˺_�"������)��5�'ܮP$��>AT� \3�iN��#�F5-���I�ʒ+Ӫ�q�qt�S�!:"k�4@����Ϊf*0�����������Td�<	�3���f�Z�˹H���������r�e+�6H�+	[���46�ڣ�2O�ʹ����M�.z\����7�Q�.G�e�^��EKHX:�A�u���~?��W:'dfh�S�±�d?���:�*��T`5[��j�%��caL0~}H��sz6oy)�� �_�d���-�����	<THn4�i^(��xz�Su���[����_�+�ٍJ)`��B�z��K|�4�����_�T`�2[��щ���am�*�B�Y��Sq�Xt<�"�����.RťW+-��&Lw������R�Vcۆ�̊�^��`�
nn�Kw��j �Âꗷ�Yl���(��I睚��B#���tH7/�F��u<��v�����8妋ƛ9�*�1���ꄍy@:�6���6Q�iD|(-���f~b`���$���8�WRy9�燞l������d���b��e:Ȝ�!�Q����#�#�ض�"O�G�E����M	W��79���R�~�X�E�kU��R�&Ǧ����˵�	2��w����G^��3�a����I���2M�Y�A�����X�X�ڶ�L'eF���t��Aм>%P��w��:�@�<�C:!f,}n4�h-y�����J!�r\w�+d�!��e�����.����uWv��a�V[��c��i!$�M�jP�?��¯��OB3
���L��:�h$T��˝qF;n:g�U�υҍ���$*Z*�=�Ci�b�z�Ґ�!��<B��R��Y�������䱶�EӠ���6�2d���] �
��g���쌫�@j��=�+�g�g�ጔ�M�4�3P괡G:i>�yVr��:�f�T@&�$�}�%̿��$�L�[�2k����qa�Y��a�p�X�7ˍtbV�[���ey�G�L]M��`�H��~e�����o������z�l�x����F[�!Cܤ�m ىtE�/1��Gp��kt����_��N�C��i��/߬���0�mr]%	/k��i1���H��,òAX#ծzs�?|}�[�|�%X��v�H��	to#BQzu���˧+'&xF��gIW��KDn[��&�E�6�by�E|f�:�����-�5O�ŇYU���9��~�(W}۶G��}o�D��T(]��.0��(B�M���-@�P~���	r��?�������I�KQ=\fᐣC��'F.�¶����x��/�(��B5x�b������h�HA�ܡ��=���n��i@U��f(��.pL5kxdA��̹3�����