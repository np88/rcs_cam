XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���I�Հ�ƆQ�FLz��IF�˲^��"��Ё�G~���
.ۤ`:�L�G{y:�0�L�x��nXY�\��qQ̠�0S\�	��f)=��fx��i���5gd�v�	��^d7�S$A�G$#���h6�nW��r�,��KZ�17���S�h��5��[�r�H{5�䥭1q6*v����8���U��Jt�U��k.u-��~ן���X1X�DciY�%x���RH��B��X)���%6�k�=WJ`%�zqz�-�,�'�i{y�"&{W"#B���4tO��Y����E��q'�-�|U��89$g�����Q}�e�{��A��28�Y����K�;�ge�ę��M��+��m�ۄB$Q�Q��ëI��H2����T�@$�mi���5�T&�,���	�ŷ��Э�ۋ[Xa,�۔�]�${��},��ik���!0*�/��К��0�����&U��L����mh)!���Sé��f$��Y�R'��}\mT[��r�o����r���J+��P��	��8�n��}-ov��/17?X�M!�8@V#0L�:��gb�D���"J�����4���c���E���VĖW�����@�?h/XKM'�"iui���!�P]�{�]�99���{��`�&
�rB|^���u���HDcG�l��l�33��^���*���7��9[������;}���捻 oͭ}�_�u:E@�ح0���j�+����?��P:�*�7��֜C4fXlxVHYEB    20bd     a50!�c�x�*X�aQ��O�5΂5�L�!�/E8L�vO��.^ᒽ�փ�,�E�}u�B�x
e���Z5I�<U�u����K9�f��$�Ҍߏ�'V&k��}����8��~�P�<�d�!����o���/������f���E�*[����KIrr�/�s�W���
h�!��s��������XS �r$���ؾ=S�hXb�D�����ᤍ�1ŀ�qg�:�Z� �c�4�v��Z��t��w���{�!����'�n+��"�fQ��\Ubuw���\�U�QP������0�mCHd�ers����d�=.�W��d��?��8�a���������N������C�o���^P,`�Ie��*��|]��qWs$<����G������0���|�e���`�Į_�x�d�;�s0*i���c)E%5��@:b.�<���*��*2Ri�<�˛����	U�DW�[�(ܓ+��F�%���!3��98�x�ڝ�*�7��*�����K����A*�Z���Ş��E*ʋ�u
�W�U��d�;���Mp�����=O) ���q��P�It�@ߐ~w-�5+���h�δ��Q�]������ R���XU#B�s�]Zy;�U%!ΰ
4p��e�b��YuU=Ā>���&#3_��lG�7�C�n��wk"l�J��7k�Ra�t������!ŵ?	�\��+��B��.��BĪR�_dF�+9�]Ծ�4.���CǺc�(*���4�Οt@k$)��M+.�����2�lp$jI��<5�p�|Sf�1���L5���|Ǒ��4�2}�4N�rkʜ��%���A�����I�p��0{���U6����!Ah�w��+�'j��%�5MW@/�0����֚1r�*̩u݆�k:T�"��ß���K�Bc�l9�J�=����Vɒ��^�&�\���W�_T�������(���8/�~�	�2@*��5�k>�b�n3g}C�XCgk���y�O{_�q�O�[fF�Ű���C��w�ݯD�ddg��W!���ʙ�0W�c����=��	Ml�� ��!��2th���z����K����]�zX�9>ũ�p��e3�e�����t�ƺ��]*C~�6_o�a��HaOK,�L"|�{c�hYb�.�N�"�m���6Yw0C>Rm�E��C��Sb��'��t � �&>l�yf�}i��x�^V(�I��x�뭀Y��5
��MƘb 
.0>b�`K)M$ƹ��{pp��ϗC�h@��C��~_N�UgX�+��O(2pdG�M��h��Y��(J���Ju�,;���� %-=vM�Ms$����2����hm�[!�	2� LW�Bʀ�+�B3k��̇��I�!<�v=�V$�jZ��]����8�c"��H?�)���d ����̅QP�G��Zc&$�N��AdKR����e�ӆ�}#�k�,r�g����5Q��O��t�����
��&����
�|��xđ��<�^׸o)��Zn�O���G�UeN�q K��g�L⭚o��.gc7Y�`�ʂz�2R��?�Q�b5���>-#ę~ *kki�p&ϊ�So1���C`���@����-w��>K%L�Wo� �Q�����Iq@@��6g�뀤Y�> ��ӵͽQ�PW���J?��Yʟ��E^Mm���Jc~�ѕЌ��|�-�H�V���HB��p�T��m�8���i�~��G��a���z̋|�r2Y��.i0�6��%�ChJ�2�Ec5�����^4�7>L�������~��H3o�[��K�YX���Y2f �z�5��
��s$9mo��: ���Wz%[TQll/���� �-���o,������&@Ľ�<#>�z �A��6\�A����12�m0�/~�C� ӴL��O�[U��p�'}s�ɖ�~��ߗ�����~+��|�Y�K�Vʎ=�U��B��#p�æ�K�%��$#@Q��T^�N�2���4Q_#T�55�����%��Y���֡4=\���oEV���m���E��C��I��&K�Vx������/��4��2$]�p_B��_�񀊘�;�LAH����Oo`+��X��{G�7	HV�%u�Q��h�H���7�X��Vfv�S�����vԤ
�}J���B�l+��bǪ|����Y��c�ϼ������ҵ\"��=E�>�����e�����FŽbW!;f�/����lWNd��߅���n@f��,v#�M8��Ճ��Y����>gޤͿSR�;L9�7~��� R�z^^�4+7ɦ�&���i5��J�hU8M��J&�w**��?2Ղ�[��<;�!<�F���<�z�&�&}'Ag	��C�K�x���D�f�)7�.�XS�O�'S���M�|X:,����a�:9����h�g��[(��Nc�� p�j�ޭ�
H��F��J��Cla�����oa3v�,���
�J��a�5���<��:����0uX>�b�7/_��](*2�X%���>�S"[b W�Y��in��G*z.���%x�أH�?����uɾ����Bp#h,�&ӆ�\�, �X��&d���B�f'� ѩ����m����S���