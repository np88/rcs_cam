XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����}�m,���sx����f�����^k���W��!�7�HJ깳s���4>���~I�C�bh�d�o˕��h9��]�2<�!���?h�#d��"~d{3`�S��Ν+����%w^X��TbD�H�u�+�Ͽ����r����&+-nt���#��#1���(��v�q��.�b��h�Tt"OFqf��DCgUOYBS������Fk�ej� ��H/c��|��h���z�e���G��%��`���JL\eM�nW���ɉ�S��*ov�n�~�!��w����g�	yBؑl��o�9��U�g���%�<F��EW��ATN'�/E"(2�w�.2Ll�/� �8I	�1� �&��?�^vҕ���G�1G�&{���h}+�E�$��)A{F��\a���z���w��d��л�g����S#^�`.�9��>E�X1O�L��n�:3�q�|jGx?���^5E��Y%S:Կ�!���J�ҽͣ`i�&�������Q��(��q�}��r����a�5d����f���M��p�Z�:ƴ_,�zVQ��2�X�3�_ǰ�~U�
�����\����K`�N>U�!Y�I������)��_���t�_���h���ϖ'7� ����<� �r1��g��Xɮ��~՚1�}�NL t��bm����嫑MEU�=P$/) +��!-�
�N�,R*�[��%H&E��V/��C�06���w�	�?
�[�uÆj'+uUk�q���-��3��NS��Fv<u�Ύ���w���Z�)XlxVHYEB    8405    1280�)#"���_��ؙ`�2�����;|�/%n�{��Y��Rtj��)�v����I���1�lW2v��1�s�JK[u��XxtK��T*����#o4��Ĭ5x,-wԿk@���Ķ4�g�C���%� {�Ae�2���N�Y���Z�-�I��*eL�<�5�����NZ���Ʈ�O�~U�@��~�3H}�w�(���F�i_Pa+Ꟊτr�{�`K�z��i�&O�N �ͼ�	<�����@f�S�">aZD�����y��߼�N�o��j��`��tT��kC��HJ7a?��1~�^�N��C(Z/�%'�nu�*��!�?bK��k�U
��G��"����J*�Դ��nJ<�
=��1�a^���Î�!���oJhqRPkg�Dg�|[��I��^�q��vp�fm��g�X�����$��*�L~˅Y؀�uf u�+�Wx֑?�{�|�Z]\���6���o�{�,� q���p?*lR�H�!����",��ж&��Js��j��"�ng�ǯ�˽H'P :�D �@�H;I���2,��/�3�T������wHp;PVe������W�����i��������"�kyk��F��ۈ9E�	;�ܛ��SgۍAx4�y8IP�f��g�T�׉F�lp����-;���-Am��tg�m^�-w^6�8Ռ��뺇�z��˱T�}З�����~����vk�"�W��-h�ĭ�CxQCc�b�Y(TE/��X��*p��P(�|���[1��(4�-�������j�hO���i�5jA����1}0 ��q�@�C�x�\��M��ډw�V��4X�'y�j {4��C�$_�a��i���b��M x�.��c��۴���N�^�jhǎI��c� 5�^�L�Υ�6d�2e��h���'������ �9���%�/v���/�8�O�  ���c�l蔝	��{��Z��9m�VD���$��Z����CM���H,؅t�q�)��b��� 卤O�0t,��gJ9dm�&���O�ٺ"���*��i6t�����4��퍶;�N���X_�q
�d)�j22�?�,�yQi�ܺ��L�:q&!zZ���>o�C���fŞ/>��q����VCd�h��0���Z�(�m��fZI��,��3�(��P�m���\��7��8���0ഀ�Qw�G�O��W������
��"X�y}0u�)�4�w���7��=R��P�)�i_�ۜd�`�A���8e�_CtS�-�Rby�dw�ؗQ8`���K6gh��ı��O����4ɵ� G���׊�xF��Xs��ks�]*�,A�ԩ�l�Vu��O1�	A���lVAui ve}5��6����h�v�ب��k:�c��Ifߩx�l�0���*��M���ĵ4����\���N�ȯ*�7�̃t>�@�?�n�����n$�M�~\�-�>9�$x9rꎢ���w�O�j�g�B��]����u8�݃ᇨ�>���ђ;?Pb7�D�G6�w�f�������B�ȹrm>3.�I[�����#!y��>�	����C���$U�l@�3���:Ȅ8�B����ߊ��fk�X2Z;����͌@vUr��#A�:��N�|fh��A�'���-��J�W���G��^g+������#;3�0�U2s}#�s#�y��뇥���-Oq3i���v�i�|�q��鏆�ď���^)T	��6^�*�Ɠ1S���E8'{�&�n�S'Bdh�!����,l��Jc�Ìӷ%1�~���Eĳ8;���5�X����O�U���~zVU^.���`�S�� ��x	a�O+�ݚ,�Ȗ�y�)f��,��Rz��K��(i�\�^{Zb"��͌?�y߸P	�[v���_$�&MM2��^���D'�W]$����9�Va�l[��$%�C�JL�k~j A
O�X�X?2�Q$��]|�c����ѳ�s�c�?��;}����C;��u��q��	�y���!1�p��\F��yƂ�UoC؏�J)�1���ێ����!����x	r�P6/�T��<A/�I�ؖ5�O'�x٪Ԫ_�ls.ۄ~�� ����1i%a1r�:E�H]/[n�!�������P(��en�ң'[~���&m=�-M����(��k�'�HF7�Y�)�s|%�7 S[��ܤ���AQ���F�Q@J�H���)��������Q��`�`�n�c�ܕs��Wߞ� :��-Cb��@��%��\R�� 
d�)�W��Ub	^��^�f���k����iDc��Z<��/��f�=�)
���3�#�s���9�d�JǦ�'�1/G�=	v�xر��Q��8$vJ3滢:h~
�(	�n��P�M�#Q�y1�\��Um}�+C������� ���r�811�d�h�2�v�#��jΞl�~�2��n�5��񈺫���=��4�ȬWF���t�J~��A�LQ.���>$���Z�20�.n�QZ`�L���� ��)�-�02���,��tZMGz}�JtVH�u�1߹�YzCz���K�q��'�iXgZ�'B�l�g�������"�(
Ը�}������R.�kX��g��،-H���[�d��eOo�x������������9��CQ�W��I<��&b�b��oU+<�Yb�J��z˨^�)�����i�H؇׏}�Clc�5�擏ќGE.�}�N@�PT1C*��7�U��{����k�ڣ�n�:� ��yO.�_�6ö�z���A�Ɵ�[��fU��:PV���s�UQ��Ɠ�8�,���� 
�LᯉZ�kC �c�o�+��SH�Y��S�kՌ�	^�/�h.�!׷�M9�9�AiO�P�me�yu��u�i���\Eâ���^��Ǻ���k	�Adŕ;}��!K�A�&�L�N�&��etb��4$ӿ<ܥ��(��e�S�W�`hnP�Ib�݀jY���+-��b���!�wX���2\o���H�ś4��?!̣��56��F�e�$mp3LBm�w��}�����`����%�9�m�}�%}���A_�tF�X�	gJL��*3��Pk��9� �s�.	�sn�%��5l}~��\�&p�d�F�������{�ڎ��1��I�]�:�/8E��	5�܅�a�lp7�n��*�W��S�ŉ���镼%T6n�����x�S�5�����%Mz�'��4��.c�D*&��=i�$�;�Ӣ�>��'�CA��M����^��0`(U��3Ɲ�z��OTOj�M:O��	�eӴ�; ���2�L��b�$=��Ħ�����#�i��A��K$�F!�Y�xc�m��Q��e]ͳ��%��Ke��9W��û�� N|�lLZ��=G9u;�����|��j.�;��0����5�F�� �W�'��H�b���m����Σ��2yS�u�y�5�*�jFq:����^��."��hS%�F0k���B��kԗ8N�!T�ƾ=1q�塇	�0����
�l]<���F:�ֹ�fw���V{6��Sx뭽Ϛ�<!)��M�&l(HCPr�m�'�;�i��j���aߨ^c�trT��i�c� �Uph�Z��8Tc��?�Xr��NJ�i�>�O(U�2r�)��/k3�d
$ܧ^�sjU�)�\��".3�d�VBg����X|�o�x0A�}dBbnl2"J6�n�;�D�
���'�� �b 0���t�	�.!^C>�k٬BFW�
���,_4N����׿�؈����(�
~�Zf�>oK3U�%�}˨���|(n�P`U��/7������}�/: ��A�Ni�2=��n�����\_�,ǮzY'Q����2z�uA��"L�8��{����Z�Y j���ҡe����l��B��Q�����ș���E9ٲ�����u�J1�"�mF�:Fp
��fE���^��r�8��w��׵Q���� ����w�<��"AD�{�Un���ㄒ2��M�;�8�E!��?0�3m�8���ֶ�L�l���W�7�b�  ҙ6����s�:IS�O�;��u����&��!��A�y�Ϻ<>ኣ�<�:<�M��y�S�>��ꀏ��k��;������BP�x��S�F�x�$��ޗ�����h�½��ߤ��|�*ǵ7�x��t��!��'#j(z~�7��=2L3O��V7Էb�p���`�0�7��!������;�3�Pz�պ�YMwK!}���Y �F�ds�̝GJ#Nz\��F(Q��?# ����_���*��d�e�r�j��^���/�ģ�j}������z�M�0�h�v5�y��?�t�_���]��G����N���B݀����^�ϥ��)[�ۥBB��r�h�j�Z� ���`�4i��ς��
�/C���*V�F$a�T���4b���x�*'�%�a���n�ivu�zթ
N��׃j'��h�=u
gB�?3��e��y�Ūɺ\�T͋��b9���$��e-��:�z�(�Ȉ�n�+�|-ڜ��P�����y6���d���k�'������$3aϫ��vV�LL$�ڸn��L��rl�t�`�u�Il��J���\yG������<N�����D��hf(���x+�:�6�G�֗g���9c�E