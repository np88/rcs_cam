XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��v�f�
)��I�4�5SXM�(|-�
�GR�r���\J#�N��^j�W�G��O+P`>����^*cZ���=n��(��#�'�lǼ���y^-� kT.;%�W�}�C�~��բy��q�k��+�O�e�ID=����E�[N��g򖚔w�}oy|1hq9����ڑ%����X��; ���v�z����h�sfCQY o+�2��Q�R'�z���J����|�A��D*D�F�ЋUJ����Ca��ɱ�q���]�8+y��"�+@�T#�2iٚ�����ʳ�F�t2u���ݢO��%�\��w!~*e��X�4r��|W��.�;���(O߻�O��A�9C��"ˍA 7%1f�ej���xy��Y�m�ܚG���x��$%�=���F�ΐ�V�1C{O�ˑ;-0��+��	��E�}ѥ�+�\܂��%�iQ�L���&P��#�����`�(������$u�)�ZM~�$�J�z�`^��ߡ��*0�|N?v٦�*�e[ᒟ�ȶ:���4�)���	�S烮7+L� gn~#�S*7�1���Uaeb�'
�QhlxEF��JR�;�O��} �,Li����Z7n���kWgp�� ����l�WO?��p�[/�v}�3e{�uGpU�+�C�ѷ&Yx@c�1/���:�Yy~-z��J��E���p_���ꪀLL��!w���~�Cm����S��겶[6i	�H����g���17����mQ�rFrD�m?h(��3���3F�y�툥XlxVHYEB    50f8    1010��Ҳ0Y?�B���x>�S����K�8®~��7C�p��W@6�E������f�<rl��@:�%|�=��]陱sn����L��c'	�cM�ٱ]��O�z��3����R9B�mZـ0����M�_-� $ȏ��#��`��#NEX}�~N�-E	��Ƭl�L~ǝ���ˤh�FK>���$���W����Y�#�����pEy2bv�)�_",�e;f0�yy�!h��v�[E�8�ՑGc{��=�G�:��X�yiD��\yu�	hX��Ǣ�g��`��<��fJ�jK�xs	zy�h7���p�L�셎�}�;K��~n�o����*̋��oJyZ��!�� ��j�ԮvCR�h%(���ISNH�V�_XaVlA����#��G����N&�����<��q��b�L�eg�n�E������>I��'}r�S��aCDqe2�]�	G��?jĭ����z�DŊ���a�e�s���j96�.����}	o�6�ۅ!@�AF�:��97r��bXu�n�����YL�P�# ٖ�Rl}畧ȃ���L+�u���������\\WS,$�9�QU�x����!��н�s���%6=;W>�	��r��h�.�=�whi��e?*lAΚU�f�����w҂i|�� �� �b��z�X��#��]HD����?UN�4Z[���TPaʾ�7�P"���s%����'߼��
ݧ2�|	�E�ĥA�,�7S|-�<�e����w@|sO�U$ar�&��@q�%����w��5d̲b}��^��Gz:=��[B� �Bbӯ�g����b�:ԉT�6Ό��x���
yZ���T�}�e.=�8���-/&��;�R�����"_��B�4��6N��Yͤ�y[`__�ʜL� i���
����P!���M����qJ���h>�c d	x
Yi���ű�Tط[�t�#0�X����NKp�x��r��X�IJ��v�	�c�?�(��EK�P�Px��2(rV�t��Na�+t����mc�vu��\�I�A^�,X�}����'�y�v�Ȭ�XW8 q��	�����+�� ].���ۆȇ�� T�'Y���"aÿ��3�p~շ�Ԫ�*�Z�`�a�	=�����p�f��SC�v���#�Sw,R>���bˀ��rva�g��R�9r�� ܤ�=���N{\n�sZ>F�͝Yf\Uz�b�J������'0���0�GX3=cO�H�B���o�aL\�l?TEqY�#mx�s�v�0ٲ��1��J�$I��?�1Z��Š�����̪݃E�ϴ�/s��	;���*��ߔy����Ȳ9N�˦FHG�z���Xq1G'*�`ǒ������2�uA�G�N���>0�ܨ�s����'-�����D �X��H�?M+a�K���C����H��M����U�vc��5%%aȷ�k^��;���&[Y�]�	�0T'C�1�\%M�O�:����y��e������~-"�-j�e�@M	ĦH�4��N��r�j6tb�������R��dyIb�cM�M��9N��J��F��� ���d�"㣂��*���1�!�Ai2��7V)����,s�(N�z���&dա�O�[�������ZZ���#�M���aS�/�GC�~u�x;��6��qO��zN].��?����CEU�Џ.�n��b�b���۹��+W�:P�]nw�N"_!�=r�H)sa��xM��P��~�2��'	�A�pE@���}Ϗl(�ġ��
�˴/�i����bh�@̢V���E��e���B�<��+K(���(ǅF���?n�Î�f�ߝ�9Q�(L�pQ��.�<{:5�K��3~�rߒ����ĳ���~�T/R�̛f䢅�z���$��3�_��nӫ�����	������5�����q�/�x#���Md�R��o�}S���e�	��,���v��� _PϬ�Gs��tZ����@-�r�M~��u<(�sK�`'!�N�>�I�P�U�Ϊ^� 1�}�'��c i�!t�j�	�pI�2,������2��f7��8�L��(P�.����qE�N�ԛ��>`[�a`4�DP-,HqPE��X�O��*�[����{���{�(�\H����� ����T�,�\g�����7�9m~�h�Nqo�(g��'_�L}٣�a�=g'ܘ}���k��V;T�q��1NP�}�=�����.��h׳I8Բ��|5"����)���Ojro�LD�[ћ.T 6�%z�Y����ʌ��<4Zv���D�c}F���u��k>�ڬ�g�k�g�ˠ ��i:8Gi��W�)h�k�V�H�B Ռև����W����Ю�<�g�9F��ׇ��Z�;�\��0��2���C*��3���|�W�F����P'��<pt�Q -�����;_�,�ר��ߙ33�����$�+��m��Rkl��J9��� >��.!�F5��Wҿ���]>��#G ,��("�E�n�"rL���t��%�(�Q\K��v�v����=A{~B��Gb^��xi��N$���E|�A���;�ʣ}c;P $�z&S�Sq����~T���&z#5���B�k��ɑ-UN,��B�G�5-��/d�v�;K���X����ݬ�F����1��#[�+��$jiQ`U�RR�ξ�S�
m�߳PjI �RFs�I�T�8��hPĵ:^�R������s��bҝ�M%q�ش3�Ò���zp�1doYy��+���%
�{�͖�<H��2��;��ʗ��:cG�%Q�./��-�p �EǾ�޼�)�!1d���]�;.
�h�S)�G84@u�!� �����wn(��m�q�s@�~�K�]P�#�s��-��0�ږv�񟌼�o7�@�$��"��A��ec��lS{y�7�GX���I��?Vi�I^�k9�~rc��R��+\`,��p��	�W�G��Z1za�+9��h�j@N>�,�é�ϴ|�k�k�tP3
w0AӺ�E��tv֪2)-��x�փ���c�Ɠ
�i�l`iqh����	�`4���[�C>z�w���j��T�j�P9���e�w䨝*���2�xX�k�d�'l^o@��ە��6����lv�����~�h���}H=��_���X����Uw�T	�p���}1^�.��v|���ϢIȉ-qwX�����C!t�h��0j�B6��Ί}���o�X���B̄������0&�/����*ϙ��W[��ھ��I=�dOb���2Px3U���Y����RV����~o+����S[�zĽ����
w�����4p��unP��#|�o���]�v�zKa��"�g�n߇&��� l�@��}��N��e&9^a�r������Fd���,����B����I�4 ��\�"r������� G�ISҥ�xi���n
�V!�+F����\=�M��)�/u�s�K<�.}��eZ�J	ޜ�	?C���}ϻb�T�"�f��;�&O���]'ǴZԪ�2�<_QU�q�ۯl�U˭]��#>k\u��l���c�KW͕4��n\d��R�d-���-rߍZ"Mm�zOU�Y�P�V���W^�{r.��#7^&�+c��L`���rܯ��[ȱp4{��=f����\���uP}����e�/��_j�9֋�e�u����r�{��d�U��H�XA�
 ���.j�X͔,��0�K��X��@? �
3���j⳻�,�,�$��8��-��P6b��*�kqn�b\y�^؊���_mp	���7���E�E6���\�H���j�p��0��$��-���.J�{0��c����� Oا��c�7K�%��<�<_��;ė�2���j�ư�����Ry$�>�� �?���٨��O�Z�^�~�Huw�Z�6����o~;-�>�i^"t�~��arL�3��\���x��w<yh�!O�p�	�m$�ě�Lb%̇�6X�8���s��/��~�r���$i��8Zkw�3��/�