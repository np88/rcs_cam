XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����+���ļF�����c��n��e<�i ߔ��n��C�^���Pn2�<�z
O�4���/���B3)\6[���Hn��Ey���h�<o"��@'�+d̐�f���N���,��J�_k.ם�Ǚ���s�ش����M7�����	��x�̱��ZǨ|����|�������fH�@~�b�]&;������\t#(A�u���S���
��$�[ȝ�u�@q����@�9.J�9�U:L������W7�UU��-='�����?��|�	�n���\Uڧ��<��u�AR;+|;��^��B��*�`l�����Q�y$f6�ױ���캵�Y�ʳ2��!�I�,_
�r�Od5d���9�_���Z��aӲ�����/�a����,��Lu��A�;w��L�m�̆��{�[|�?o�90X >>D5Z�0�}'�ݾ�oƌw��,wˣyW�E�#u� �q5��YmM��	�7"�U5y�ӵX4g��O�Q�!c!O'��2),rҽv^-��g�2�@m@\��f����!Q�����B��wq�cU�����N���E]�ዔp\�j8���iT�������/N��b{�{qm4�Q��J��G�7�l9D!n��^Ǻ�eQ��;1�	�+�jr ��r�,���g�g~B�BVd���Y�N��!f�Y�y|��bD�h7H�V�ܮĎ�?4�f�8�2"��J!�::>G�s�{��R��re�v{�;���id���W}zF��"�	�
�T�05mXlxVHYEB    9732    14d0�s��k�4Q,p�Gq�Fw�z�9�)�_v~��[qP����'u���a�
5�n�O*�K���d|�6���>�w%r��	�;P�a����\����a�]�� ůS��<����`ԕs��6?�o�U�<���e_쁠B�0_�GU���*`�>R�(o�n�������M�1Q�A#��)�;����ei7����c��9�%�4[�̺�<�f��u�S�y���ܵ��ӆ�E\Op��o��!��5�s���2��8�
�i"Z�l�Ґz^=���Iq���o���{Go+H,���0a�H���W��a��Y-�>J�I`<�Dq��Qg2��)��G@7��@k�2����Xy_����^+s> =�?3/\�#pJRȾb-��I�ߐc���W�Ll�1ǵ�|X�l�B��H�����TshY����⊙�'ǔD���SC�.=�`��T���>Uy9��V �#n����%�҇~��3-łձj0���V�h�
�;�c�Ǜ�Zb0�1@��=Fx�U��z���[���5j=��:`G��fjZ�S�(ˆ94<1��e�@g��x�	�l�S9i7���Q2��)	~�x��L��ԤH�@rP̷�xQ��|H�YT�!k��"0eM��%���p�.i�Jn�eB0q�M��f�N���2)�_֪J��z�=E�[9#ݓG0����:�J����qmM�OM�)qڨqe�Д�s�.�鸢u�������Z��T��=� td eV<���)�]Px%|��:?�����Q�n�r�������Y��0�DL4���8�.���]eo}~�FE�e�r]L�O��p\���^�5}�	l
��3����A��n������U�D A��qJ���'"'o�C�Ć^�_q����r�CV�<�K*ϣ=A��a�U�[yߨG1G`��m�WɡY4��էM�&�Y���|1_��|x&]p"�� ���~�U�-BݥC{��	|8"X��l�欱=y�%�u�i~MsԠhKd4�6�Ƃ�cE�aj�/���b���Jt|�N+��>O+��"��~ �P�"B���{����?��L���+�+����2.�}`��Ьm9Gz�����0�;dJ�_��;�n�1F�B±���L��c�Cu{w��t�����/�I��AD k��P���dZ^��
�����V��X�uƅ�������e�	�����pL-e�"���r�&WJ`�zʁ��]�q
���sֈE��Q,�+�?�J�ē�\J1s�c�P|���^c�~S�Le{#&����h
�+ɋ��V{�>G��R��V~Nb��*Q��b��:�S�z$��iЧ�w~Z�|�)~Oy�:�+L����Z�"E�x�%�%�,��j�R)�z��P�$l(��	*��ʾfCi��(�(r��j�jq	������D�I4���2�A+k� ��)��?(T�\�
��>Gvm��Q���3�Rnς%�A�/R)6 ����Ps�TF	��}-]�U��wK
�IO��}�%��%r*�@�%u�x�`>����g����Q��6��qV	��}�ڎA�֯����z_n�|�����ҷ6s�ml���a�t�����MX��e��a���3$��T�;wC��,�k,�K��J��������5�jr�W�}�%�)|FP�J�S�痖e��>�pn����YNwiJ�de���Z�7���n	�	���pX���	�Lma�_���8�����B��9+�eܽw����zz~`:ZV�1�5��.��tkd�fv�����$��"M����W�H����r$��S{����)��N�n]�pϲ��~�3+T<��B���vpEH	<����v��� 0�&/�\��т�WnVt��(T�D<�
+�}�b����Ξ��$�[��vܣE�8�m���}�M~[L}��s�v5�����1x�;a �
-�艢�@v0��j-������#:ZH��I��y�hk�	.4���s������UJ_P����&���?v��mɃ��Oҵ8����>��{
�[�X��_�^L+=_/Y)�&�g��Y޹|���[�E�ާ��Ƥ[ ���p����������7�7FŁ�p�q��%�a5�Q3��Wc�+�_/�ށq�iJ�����Zz�^�����
�D[�v�ěi�P�5,8�����".ZP�����@ǹ-\�y>���Dxֶ�WZ;���{�5L�Tڳ�:�C��g��9:��j��GI�pRl��/h�V4M�B�t^(��؎���RH�;"���i�w'�~�P]����i�a��� �jU#��&���n�D7��=����AY���A:0��$���?�%�B�5m��_������l�K�fo#s�s�1�
f'�G���"��U�jt��z
<�l�gT�.��K�8�j��XMH���C����0�r���e`!~n��ν��/�^���i��@hW�Mj��<�6��T=�Bb�w}x��e*�RU���\K���;���h�_��Nfq�^�z�!ґ��
w�+[����e
��o��=G�2�- ��}�8H���G1��Cfԑ_��TәfP��Oa�h�<A4��������$���-	ݵ'���r�$R�y������h�h�q"#d���̕�yv찂s�(J����X;i7��t7����`�Y�����k	���W�ά�p��ɥ�t�%;�ҍT��\�s��t�s�
:"�Kx�+Q�:�5A�����#���"��E��}\��.#�Vl�p��\=���Tr�:Ӽ(H\q߁�-hX_%x��o�I� �h
��B�}���rV�#T�'ӄ����"����P��y��H
%�d��q;��M���-P��my\�ׂq����)0 }���+[�����,�����u�È^��/�u���X��ν�<�0��><a��p����r��n�;T���tA�1�|��ǚ%<�uC#�Ꮯ �V?��M�s�J6źe���kLi.3�a;���4f���#����������Ц�r(����6���(R���+�)�������$wG�;�F��w/��-�>(����^����� ���^`%����Q� (
�WNo�gщ)W@�F>ؗ�����\d�A6o_�E��9k����i��Khb��h6�Jޱ"�@�Y'T�P��S����sX�q�D�.l��p�������ѩFUxi�]Z��e�_�����%c���A�0���|?�.XxC7���o�P�K��=55�nY�����Z\���֣���l�?�k�'���O��x�H��ɇ��y���Gp:0?א�T���+�9"���O{���Z��"Z��>�I}�|:Ѥ�x ރ�f��球O���$���X6��ȍ��!�Q��~,	N֒�b�V�Ε1\|6�(�YKc@�}��6=01<�8��QҦ�mywN_?KĐm2W)�l9���ZB�e��$�uc�R0��}�l"�`�A?eO.�;�k�;ʹK~��{��&���7�`�c{;�P��Bt��H��������/�P55L�xs�}�� �W�� ﲔPB�
u�JÇ�a�����v7�f^�R���S�dq�@yL`%2�����w��X�{y[S�NoO�g0(B̫CM��-݇7ó��2��0�0�3d0� %>��]�s�@.���)Du�w�˞�~��~���r�X�_�����L����#(+�m�3�+�\-Wzy�|�D $���$P#�w<��#He6;A��X _ű�j�&y�����ٚ,��52���.�v�Dn���e�Tq��p~��]d^n�
Q���"��U%͢Qs&Y�Q�÷��xT3�+�xT%���'���/·��N��F|n�J mլ1Å*��07m�n�9$�Ӯv���I@��(n��W��C���\O�!�~f�ƴ>�p��n�)'ewⱨ���ӎ��w^�:�,}[^���ɚ����*�<���l�]P��l�[9m��GE�VE���V�Nbq�N��T��M`5�oi�{U��������id��o����Ș#��U�2��&��6X|u����=6��P�c�>�%���L�m�1c�n2N����'��~��2ĉ'm|���i0���;;{�P�0L���Ȱ��#�ET\W~%�ܪf��ˍ����[�&�Q���t�������?Љ����(� �z��(k�s�����̯���o�è���9KwY��������o\w m�9K����C�nI������ԇ�,Y�%�%�TV���y#%�Z.s�.@��(Ai���;��YU�x�v���"VC�U �(��]�٩x�w+tx*S�n?�o,u gG��&�)����̥�A$7I���Ya8uԲ����Tr��Z\>�N�4��^�زeG�_{�Μ���A�T`��ߩҞ�h�k	���֜�C��$cF۹_�&)��tn,H�6$6�9'���x�^�hjԔȚsv��	 ��b�TTcDɀ��
���ǹonP)�Fy�����"~Y���B��ɶ1m莻gd뚵$� .	��$� ���k&g�oBK|�����������P��h2@Y�-�����;��a*FF������o{��-i		칻�萬H�� ��Ev=ld��)�eO?~�f�:就D#�X�)��D�p�޻%��%�A��eh���_`�@���%[�Q��U���y����?�мO���v�K����cn�{�6W��i�0�h�"gps��w�p��M�L ;���(zq�-�@_c2�@��0�}��SQ�����[�^|.�Q,i$܁TP��1��<����@:�{g�J{��)r� �؁�c��b��{��n}%�o��Q�c�T������<d�[�H�lOZU0te������K�d
$>�%���LE���X�P���<l��뢇`9��@]�f�5�u�~f�0��1Zѯ�mZ������F"TmD��|�e��^��8K�e��3�5�+C�@aL�ɞd�Zo�9�����L\�vI���U�&�A�0��֝��~C���bχ���PB�q�x2<7������ ?�ѥ$˖tk�>�f���,lW��Jl��EV����q	�t�'Tg4�l��E�ŀ��*Sd�iƶq��� �Հy��n&��'�q�W���Eq{�`��m6�c�US3,��l�w�/��M�Ԝ>Zɣ���T7{D��R�
��