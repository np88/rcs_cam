XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��~{�:凂At)�#�3��oA6�'�2O�����!M��hpX��!z��$���C�iW;�5���'��r�ܿĖ;�b
t0�0��NS~�\��W:\F�� �}�/��&�m�+�&<v�6#�WOGA�#��&�U�ܪ�C��@Y���;$������sH�dlU�F5�m=��d<X"#��n��n_���Pޖ�ؔ-�Om��r*�D�Ő���V� ��5��<2b<�4{*����Y�vH/7rW��3a�9�fV�5��||�f����E`[�C�W���y̑�w;-Q��כs|�j�?���{�BlZ���_�I8�OEd�ѫ�b%=`�t�a�wv1Z�0-��>M�sJG�W5�	�y}�C��W�|]�A��y|�-��EJZ.��:X�&g��-W��/��rU,P�x�Ė]��Y+�+�N��֎$9�s���*�����?ʽ��J�*9�
&�$�MeʦP��ԚG7�|07�9����z�s'�Z9S/+���<�$���Z��g�õR���Si<(We�<0��=лt)�U��D�d�r(��!m�Њ�j֥��;E4�D�$���'JIG�3Ok�52�2���J�=F�aqF|��"Ⅎ�t{ �s�!?���ToE!���Ϗ�EBzi��v]6�l�s����#�__`dDU'H����q��<�SRW��z�U�0g���5T� �IQGN�Y�<���0�iz�M��N��9j�-.�C�\����d�O�u)XlxVHYEB    1aef     950�~r`��V������4ЁQ�T����=Ѓ8������[��o��q���&cg\0	ڕ����l�3�}o�`�0��� ^t{~(K��w�f���ANZvI������M�������,O����}�X��&w2T��8��%�Ҿ���C�X�|QZ��{���q��
��kn����Q<±~T ����yw<3�̯#�`֖����6Y6�-�Zp�M��ی~�TO�UM'��CxeȜ�X���eL�,!����T�1'���&����n�>��-/����ި�o��*_#��i�hb�T�hQ�y.�=�� ��T�
�E|��!�\m���Z�����͚��/�ū�nL�W�W��`�
�r��k�E)9P`!�� ��N��~6��H���1L�yq�5���٩��|�T�N{���dE)���!t"+M�"�FZѴ��a�>�',u�z��J4ߏ%S�Ff����K���1�~�E��#a/!���nဇ9u~�;�E�2!�RI�����W�U7�骄��-��xZ��d	s^[��22Izk���&TE��ޭ���0D*���8h`Ja�O^6/�囿Iȶ�-�18���Q�m7d�%�-���?�d䘌�~�N��~�_��,A:�2�� �=�t�^��8^y �Aݷ����;�n�W0P4�`?���T�_�PJzH��g��R@�C[b�Za��o���1F�O�4$��L�vt.F�!k9T����(�ϩ�˨�/$�H�ȸ=F���O��{ +����aM)�y���Z��h���P)�iӋm����րqa���a0`8���娌@�s:t�f�-T�)�[N��Mݖ�r��a#*�!���]�u�]e���8����#�3�W?_8<M�(6q�N��1lOWPi���K�{��i�!q3�*�I����/�;��Q7���Z�����������$����:l$[o �v�aX򽌢
���G����s���L���MU�{�JC��{� a�H��s���,��D����E΢�vņRo#L�,�$G5�2��β&:��bvb�����z�1��K��<�:R�=鰊w���\���J�n��`��ג��ma��`�),�o����o(bk�)���X�M�����1��^(���92h�z�Bx�fԪ 4�3h׎��ֹ�K,��z��9�&��;r'�;p����B<bS02?hb�x�.��l)����E�X�k�+,밪:�e��rH�c(:u�/��A�¸C�y;y��;<��3��L7J���n�����ʇ<�U8O����z"��t�5�L�t��9Gw���A�3�y$�v��1![�2:��H�Հ�aB)�쨕���"fQ��g?�h��\�F�sD�O6�wgI�u�os
�_8�1Q�B� 	'��zlW�>c!vcò��� nzʤڸ3@	�ד�ۆ�?J�����{�p��z�Y�E��W�}�mN�����ntfY����U���[�I�6���x�M�y*<�u1�,�LC]�@�*�](-b��x�M 3�Td�|R�a�b=�B��<�SI�}�5h��@ Wʨ:��Fj�k�Y�ߋ?��
��cQ2U*�~�׌W�����b�j�C��R&���З�bx��ߗѦ:���c`�s�6�	�l�^�M1�gPʹp}�������M[��9��v�<������y��cz�^�J/� �ǽ�����K2'.�n������pnF/�'��!r}~@O��p�R��v����H,����w�N���}��,/�j�t��������W���p�����rv�(����[Px�ZL��z�nL��o���w|���%�O�Z��0AF�8o�59������CKr��� 0ȜUuo����Biy�\Pڱ�@���Շ�����nq���\��T�b�ɣȿ��?Ԧ�tuV�[��%��!0�\�,gnF��h?S#W�7dq8�䞲�1S"�WB>� ]v#9����_�2��J��v��� �P~�o�* ��/P�v�6r+�ǉ*��t������i*�����ۻ�U�٥�-�i'#\m˧^Q�&�Y�i�f?L�ަ )�t@!ϸ����r�2��V�g��\S�?�����՟q���)ADAoC� �F���+І�}�4A�I�2�2��Yퟦ��w���u.��,ҷ���䋲jU��B7��SP �ݮ�S���>S�)1�A��-��)�	��vFþ���.����KƔws�a�6b������޲wܲ�`Q����zVr{� �c��"p�u�N�P��x�j1ˆ�i�a_�W�J#���f�W�fJ,�\�Q"~�*��䑨�Ix�բ��$�~