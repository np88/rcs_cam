XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��B�dXp�[��窚H��R�Ȍ��j�/ʝ������i�>W�x�f�X4%sm�ݼ�D|����Ԗ0���m�\����B�7����*2�Zԣ�a�Z۵W��ć�b�*�E��J^i��[.p�u�X1l�䨯�X0���q����B��(�2����%��hTҵzn*�.X:{�?�r���+�)&"��X=�ٵ��SՏ�D@T��!�/j��.�2{��Na���a�4_��������kFCE`!R�pfj}��1"(��O&ߦ�ԏ���5R�Μ�|�,`�o׻������QF`���8�����A�E�G��(o�}��9�s!�)��X4f�,���'�M��8�E������;;)����5vez��<�fU���&�R֋�E7Xe���R���F���{F�mf]��C����dY9�M��������I�G�Fdܗ&"8�������&[rj&� ���IG,l�`�).�MJd�"I���v{U�s�9�w� �.=�d��-bro��м�#.1�l�z�c"��bA"}<����_�cmڀ
/;06XY��#���cՂD9#.�1���x�r�`^_�I�����`������<��������9����`�]z"m������?��j��O(<XT��T��l�|+��ztH�|��nn
�ҞX�dS��e[�k�>�8 4�|�d�-}��=�^��U����ږS�y��8��n�gߘd��ؽ�67�q���2�w��lȪ<v]XlxVHYEB    1e9e     910�(l4��r�a�2na!U�%�^�H�r)P߅t%��v��84R�YeQ+�V���9��%T �+��LB��:�ad ����S�̙��ʕ�xn��B�=�2�_���6d���V��8scE{��~#���h��pb�	��Q����G���]����t�QkyH�=,y+���/�a)��z°��*Mw�����"$XOe��O��V܄Ƥ�q\�,vj�V(�-�YTeL����"�J��,A���e�O8!�yv������C0?���A�\*���k`�R7��x��Cs����u� ����6�TD��@|�~�ھ9�<�i��+qT�wtl��a�\6d:w��'tt��/Q���^��B��e����F�MTt�5$�<�����g�r��qIq�����J))\ʥ�B8K�Jje)��b�O�$��X�X�����:�c��s��򦤙�~\�`a����4ᤞM{lk��,��W�H���3��ɃNx��=��d`4
��`JL%�JG�xM
P&o���:q���e��@6���C�yC��+�dӖ2�?g	���>��V8����=4�����1��$�*= ����.sp�,sm�!C�s�{ܣ�S�џTy��Qf"ֱR��X�M�q���m��f���1]�B��~���yz{"R����W�7��P��+4)�ዲ�!�P�+^�I#9�aMo�s���U���An [�6�_���* �Nr������Ǽ��r.���H���F�������|�bv���_Ũ@�Y*B@��ܨM�)��G&��?Vl^6.Q�OIhǝz3ֈ`�a���I�	c,�"2�+5��:��p\U5*��O�4��������(��b�JJ����Z��Up��W,[�.4�q8v�?Ld�d��~,Q� �L�W�Ѥ�,'�Q�x�%��5�C��]��k�ň���G�sqm�L"��wz�V7������B�8����eN�%��;�T`e&uD�Z��&��ǁ��#OL����an��O�@k�RlS�Z_#W)�l.׭��"��g�)���x���Β�j}����?�gSmѾ��l=��Ӟ��ͨ��>%��q��'y��os�a����KwNT��߀���a�2C=;d��6T����t.Q)L�*�}�-D�)�wٸ)�U�"�J%��/F|Q��14Y;������2-G���Y��>�D�����Pl4Ί��Zsl�����.��;�~�ehr"V��9��LS�a��¢���5]LgV�U|l5������R�`����=B�f�"�BH~��X�w����O�[I�9��~�&�r�-�pv 8$�:
GA�4�n"�u�����s��Kq�7:}ѹ�b�j-=f��n�^&��L��ej�Q�E���y�9����E�0%�9��Ѝ���Y&��_|���w�'00��ߏI~h���e�#�r	BB��dB d��j���u]�)?����@.*��R�V���ğ@(��+�����e:��E*3�߶'H	-',u��ȲHaUr�Y�e'@?騠��}�ェ�|��֫�r�p��%�'-)J(E��30qP�3�˽ɓ���U�Ô/EM�)H�
k�%�w�b�MČ�P�p��=%< �ܑ.\��us�&%G�*2���?���bq��Nή�.Q8I���b�Qh�;��>�2+�{�ؘ|�Q�3���)?}Tp����"/ye#@�8;�D��u+�XY�<�3�u��^镵��.������P���l����I���?�p�(���=
��w�F��G���.ʸ���kb�c�@#=��\����9վ ����V�iIJ\{��CM�B��w�����o"����l����#����3ȧ�e�QXw�̤��r��o��<]�lMv_\Jɴ�J�I�u�`����\1mkN79 	V#e`��#{��3�>���
��1�븜���*��P)�'���[k��1oI>A(�?i'aa3�c�1��peQVz�IiE���t~"Jr�a��c���}�������~O�q�h,�|��|���3��8.�G)$�� �r���}3hx￨�ji2��`��k\b{1��j�����b���{K�D�����s)@�)��w�Cl�6��X��<D�)�R�1�A[($r��z*�{�S� c�fAd�2�������~��j��F�t�ɥ/��W�Q���H�BaN�F~�=�������&z�����j��m �k�x�M��R�Fۓ*�V~&�oJ,��B}m.�ʩ�\��AdgC����/�X��