XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����.����u'%rV4G���]���	��-�xX���X�v�^?
�G�����/MI�MtY�H���U�� �_�m� :�����0=��ǌ�	=u�.K���)��:�S�U��x�h���?���b��Ů��Ժ�F�l� ���d~�-���=�������y�z��q��.u��|�I*kC�W�S ��<�Xw7�3�7X�)�.�gQ��qS��N�m	^Y1
=/Vx������f>�Y��m#r����� � ֻ��1'9=0v�6����75T�؉�����ik@2+��&�f��ؔ,Wﭦt�v�{������i�����y&q�~�k�4XQr��4�Af�{��s�Ymd��H%�nx��* �i����S~c�\l���a`�L.�bW%�[��ab�I|G�y�G���WCSV��8�,z��ʞ��+�28��;�E��mz�=\��Y��ʢ�/X�fo�.��5�CeD����K�K_V���4JekݤVPT7��c?qD�6�ˬ������e��\���+�Jic�b�j�^��f#�@t�\Y�h�8F.e7'�\��p��p<T]g�O��f}R2�l�)����0�(�؄�7�������n��ח �_��a���7�	���r�Cwq��n^�t���E�3�k��淠#e��Ф���k�"��ĔrP�I
=�K�����y�?*Ϭ:�}뢙�a^|0o��Y�J%}D��ѩB�x��t ę���C�B �s��H���XlxVHYEB    5694    1280IO��ZM�R��&^�/o4-�s'��L
a���u@#'Fǘ:|*�<�I�QO4
+)�n����a�lX�A�҈�u��uJ2M方r֭nʹᄕ�2�f7��#xR�nڮtZ%@���8s�O˱�t����[o�&rDGa�<r*�7�6�����(@HҮR��|�5O��>߾{���$l�t���N�m�Z/�u�����%�lc�@�owɂ f�:H3�뙄�az�eJ�6j��p}J��܅ܕ��/��<[.m(�l��Y��Vm��d�& |CSߙm�LV���:��uM=TK��(5�3'� ��JP��ΌL�Q��<����1����*���2N�M��1�9&�������ˏ����b�+�Jgڳ������x
��$i�fݚA��(���v�Su^&�Pz�S���}��m����C�-�sP�/�렔fR��d������i��䡙�2�j�0
}]y�b�b>�e�$�^��;���[O�a�/ژHf� �����������L�@�����y'�,$Eג���TT0�+��EW�E}/�R[ wM=����*���0Q�Џ�{E��'�g����]:u#%L��c��B��z�!�l��9A_�S� �-MWb���WL�E�W���Y�z넪�(���[I�+�����~�m�]�e�8_����Y�DjB��.���D��ߟT�
=�E����O<lNi �C��t�o	�o2��7�bj�����}l��WI1�F0�O� ��E�8��zr���X��P*��M- �Q�ᨡ��oV��������G�"P�r�xiOt?�j��@}+	�Yd�isEo6��FBϑ�����-��x�I�%D$�t�F�z�
�Y}��޶6b��9Z�c��
Ym���>-��d�_�?kSϝ����E0��N�Y���1��'F�I���PΗ;�(���$~a��������۰�$�eg��h=����y�����⻏���rs1A>M��& U�Mҙ��n��Òd��	�_DE��j�p�.�|�^�)"�+��iCZ7���>���R�F�R�n���C�(���ؽ3ʱ�M�E�����k)bH5&�m����No2���o��k2���AANao�%��{]���P�G~x����H"��ɇ��wP�������G]aM�b$T�nX�����?��Ӂ�.֕V犝y���D�\:]M���³jЂY���	�YQi�܎��A����~���%i̶�k�؅���yZ����睘p��_[�l���Տzȍ�T�M7�q�@�@�iZE��y����+����]�8ӂ�R�dޅ#|=M[
Ol����U14Y5���k?�}bw7-�����O��a���0+]J�4�u�X�L����Ծ�!�}�#����;�E̋���3��es�n#$B���}��di5��ru�M���G���p�nɓN}K�'���^?�~�%�M��yQ-��4(��)���l�U-�u���i��=�E��� wߺ�_�������tܗ���ғ��m��v��Q��_�`Ԭ�U��tT��d�j��O�����iNU�֦A�YD��9ڪէj��c�ϐ�u;���?n�t�9�&�l���F���x6WY"��E1�'�bxٮ�ݐX�5%���@�"�n�����59W��f2+àd��p���[vT0�+Èi+����r�Ȧ0g�Ur{�EG��ڋ��b�D�h��];�F�k�#D#�	I]SA�n�]S�F׽�>]ٚ~�	�1fl��OR����ěu"2A��˰����{l~>%Â��.���2�7n������b���8s���j&���itV}�"�*U�������XYg?�i��oNG*��|抭j"a���>�E�s�$o9:u�~�9�	Y �/L\Eg�gF�g[��C����Q,̒be�YR苯6������	�>y9����h���p�ⅿ��`T�)"�|�ͫ�dd:	��S=N���I���0��w,:�5���\fN�BV��7��i.�1�˪;4;\S��Y%���.�J�J�p����K��&HG�X]۷��I9�s�ln��Y�k�P!�f0����,j��-���R�܄W�ыi�؉�M�j�H�[k/��=˅�x������j!�,�f�9j?�v �>�u1��淚m��-�����h��6�F`�'QK�v?�i&�Ya6|9�W�=���z{Ңnn�u�k��'���'�x���N@�&�G��6�в�!Ћ8l3�����8�}��=��j�=��;�΃��_q��M����Mn�D����Fq�"K�%4�Fea�2�"������4�<�%we����=H�A����o�FnIB�����a�*�F'V�h�oRBr.�z���#/v7��1x,���z�`\w6S8�=��%)���*�1Ջێ���<���KϺ����I���I
�]Hփ�G��� t2
�=��L ,�]��V���@�×��3f��i��U�����L�5��2�v�Nt�>{Nrw1�y��:����n����+����W�e��ȾC�hn�3K��ZmǴq�
+��ə������ �ۨ�	ZJ�c�7'�����=y`h�Vi��k�vUSїQK����l���C��{�0݈��F�K6hɿJ]�E��(Fh$�S�t��8�vӣ>ˌ���6�s>y�Sp���c��
	��=�|�E]{���H�-�5N���'�� ]����Z�ʹd8��b��Jv�H|r&z�#�w���!�\�U~�%>�ªc\�^��&c���(O�Y;<<*ڤE����u �$g]6 �;�� ��]��	����C2�
�QR�n�o�@a�>U���
K�&��Efؠ�V�}��1j��+��3�
|��l��M%(�6TV���(p`q��m3�:3~�F�p� $rLXp+��U���>�J�넻EQ������}pɌ8D�Ak��ha�P���	e=[����������g��>y�:ɐ��;�dJ�T*	ǿl�^�UO��13��/�g���ܗ�s>%�B�X��X�쉇���x~N.Iu���ӶN���=���K�R��ݥ�aHYʷ0q�jU׹�6��S4�g��� ���o�?t�)R�7�R!�Ai�3�7Q-17�`���v$�LB���(ck1���a��/q[��-Ϙ�m�S��u*x�c	^F�����0J	O�֜;Jo}���Oj�K/�sH�SB�70Hz�V���s���sV�̖�4_)1��&:>��][���rw��!V�?Ka��ٌ�P��4��'^��	��!tl�3�u>�Ȳ#��"m���ײ&c&��6�]n�De�Y��)(TR�~5z� ^u%?�g!�Ϸ�K.�}��8�^F��V�5�߳�Ǩ�h��g��]Q@����Ҵϥ�� *�jU�� |q�F��k\��e�q�G.U#௧d�c���� H�^��D�6o�_�ݱ�����lCj<��b%6�XfF'�l=4��\@x��[Oׁ�����#K�b����Z1��W��}��2�$���5���F���{�E&�Nq�� ǮX�/m l��ʋ�k=ԝ�6��q$J���-B�0�(R�����Y#׆o�J�㺍9l
���%����s�Wh�+��������P#�n���)l��M<�0X:�v|�c�Y`�qb���g��,'j��m�ڷ�QP�7��A�4
�ޜkg���c��b�E����RPM[�Ձ��D�凝U��xTB��֍0� ��,r���jV��q
xd�Ϝѯ���iТ�xaP��K`W�ꜣ��� �\�OQ�{WÿR�r�Td��Q�:s�Y���P1�?|�׹�AM�n0[gkB��5���#�G`����_yJ��b�O%,���u��߈�/"�3�{y��>�X��/)�r�q��~�9�` �o�������n}��8�9H�/zړ�8�ۨ)��u��M|���>	���]���Ò	�ԥ�Ֆ�Y��O\n/Є<=��z�\%|�B�#���۴͉�z���x3��&��	��PDBW�x��z�z!Щ
dp߬�S���:5�=��ز��_�[.ې+b]�����6�����Y
�M.\� �V�c����5�h��n�R������c�A5ƴ���E�� �tf������R�}K�Q�,��E��_'A�D���\h�^	����� ���:��I���ّW�bצ�s?�\Z�ٜڍ�}.�w�}KhQj<2�n��`�ނC��x�㯇
�Uv�%�(e� 4W<J���]���<9���R��]=D5��?�M2���׮.M�돪0a��>��G��D֥�ɎX䮔�㡑��_�T���;|:ax��w]2�����)�Ҙ:�b�Bo�SY
:�U��~��H�3�	��aX�<a�<��a�;��]'9Q9�D�tR�uִ��QlF���\U��;�;b�uY���|�;��Ğ6���n�,��L7��\���[�s3�.C��F�`��V��k��h������?���F��#F�:�ijA)i;���O�cU�1�,'�>��jC�FT�� _��I�+���v�x�LiI��-΀^����۟���on�LS9����Y'�B>a,؟��Z:����Y"�T0��