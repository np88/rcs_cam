XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���ܺ�N�@@�4i���KvR4}����z��1��q8Z��Y(�R�H���dP�2����}K~�8��o�8���ᶬu�,:�Isrz��ܧ�wq�j%�zQ.ol�:J����`�P�B�Q�jny�5Q�O<�Q�U����M��)�I�T�b DZZ��e��j�b��<w"I>�,^��	+����­|RL>��#�v�*���V��fՔ��cmD�Y�DR0�l��~{�����7τQ��	��z%�����8iU��y @Ô����q��v sa𢍪Sˁ"1rr+A��hX�ſqK�3r�pb*�I��GK9�ǻh�J�7��� �t�ռ����X����]ʇm�d.�������=6=����Ԑ�>;��޵6m�~�K�ٍq_-�!��
.0�*L��f�� ��f_�a�vUqOG��>*���b���h�7$��W��xۣh��_��������΍�i����`}riaD��AaZ���TxH�E��5�����Q���[��]p`ҹ�P�hK�R���
�Ip<�2u��*��0+��)эPw�#��������� �gks�$F]c�����)����2Vѱ3	nr7�LJh_%�$�]���a���m95t/ƬTg�O��ʥ�+z��A[�8G_Ԛ4���M�p��l��rfc��_4��PW�DC���d��휔l>����h⡴@(��� ԅi��1�`�^lx�i�ʎ��SgN^u��2_Ic���a XlxVHYEB    aa31    1e40�ǡ`n|�U�<�?H�b�<JA�wIݺs����xNe�/\ǳ|���V��H+bػs��q��e��Z����'"N"jg��ꢳ�c�C�N��o��h����L�$�Z������@��z��e���1��x��~<[E���>2�#�W�4����sT�%Q=���q��� ������� o�@A1�"���������93L��;��^v�mطǭ�M���t�$<A�΀�F��3��
��""x�m������F�ϡ���ऀ(���j�tJ���c�@��6n:�����mn�aǦ�^Q���˸/۠�p��X���"�~c��`��-Ԑ^¯���ĎOd�������'����RG���*qg��x�K
�kr��	a�uZb���h��?&sƵ\k�N�c_0�kw��-����Do3��+�͖�W,y7�W3iC?y!Y�����KMT�����܊��ʘݑq���=O*�|�Ky�9oi!����KI�����w!�[�p��✝A��14�=�'!6��kg�a-���J;N���Z^��ʻ��B"����$����c�^Kc��&XMv��=���cֺ5	��tu�(�y�;LI�ݨ?���|&֎�����X�Y�Ħ�e���(��X�d ����6�F|TF�+'�=Ga�[lK5�#�Egf��8DI@h[l�2)���&�'�*�m�����E����}Z�3m��N����hU�S,�R���c(SKch��_���1�ߎ6L���xU�=9q����T#s@�6��=�,i�^:�����!zv��4�_��V���[�{�8�e�t��j�Q���Ȯ�k(���j��������П�$It����ĉj����p]�u��c�n{�h�"K�}!�6�m�����n�D�5mf��aK�f�� �t��l��e��B��֥Y�Go�ڥ����`7���|J�j��`\�tEo�2�ʱ�)��X<�$�q�8YiL��[����/kڙ�¼�㫀�"4^��w�`�=ֲ�?�&�r�p���V R�7��������Ol4m���!�@���J�+��4)j�~Wtg��ַ��]k���� ���'����E�^��7C�Z)�h���;�B}	N�v\�������z�K�2��9���01<�1-�N�ş�*d�ߛ��Q"�Թȧ?˼S�p��.M��L�ː!�n�$,����D-��jJ	�R+��b@���};~4#��@�Ci�C�jY���:{⼿>p�4����R���7;�۸Y6�~�~� ��b�h�� Ɗx_,L�Z0���H{��1���錒P�D�X�"����Bl�z_=`x��o�/[�?�kF3ea�Ϋ!���=�U|[v;oI0O�f�-y[d����Vf����%�VS]]C�!�*ik�MS���` �ͥJ���
�.�_�,���0w2d�C�k���	A 0U�Sh\d/�'3�pѽD����l
H�[����������*ǐ��K(��I��>葘�&8�CA�Rp��C��9d
^�?hi���o��o�-8T�E�q����<��|]+GA�Q���U@?ŕI��Z\�=x4���M���C��2ܩ����Y�5��΍�5ZiB�� �rƊ���z�M04���h{�(r��rh�]v�ٌc=G�"K[��I����yn���C�7e�=�O��#����9��F�	�m����������C^Y�"����8�yG�/�σk��ѽ���@��DJsp�f�bPW	�ci4��݃��ܠ��QD��l��%�S���k�z1��C�A�B�n�I¸�gZVp�;�lϝ�l)�w{�>�~n>id���^n��{p3l_4�@a4D�Ә�6	�hN��A$F�����N<[%S���T�?瓚t����ih�k��W��J�$�Z�aὶ�y-~y�	#sꤋ��">/�)O��$7S�>����������x7T9`^�2��>Z�2
ِ��ø�Á�'e�j���5��������n<.�����|�)�׳�t����?v����x΃ۇ+ܵ��.��mn����&_Pk+FE�����y����=h�m�	����	�.')���$JUVp�R� �BE偲����P��k���z]@*��E�I��l�&;x�x��2�4q+�e���p ��x֫�Tx��Z�[���G� ��_o�HR�:j�mw"�e(�oZ� �Ec��}�F��mc?L�c�ڡ�̒/:$�V5����I8u�����8�S@���px��I�jOHh\x�=�:ʝ��S_b�z��:IZ�HsV"���3c�����9�e�����a�d�B�2�*C�$ʳ]gG+BM�B�B{�D,�я�S���BZcKwc��D�ʼf���9Mt�*+�$ء��`|o"��v^ё��4p�p��b��S� _���;�e�¯�G7Bv`(f����T�i���4,�9�����F%W��\�%�b��z�C4crE[���rD�S����q�U�N��!��[@������?맑K,ݐ��
� �p��`�Y���e_����G��a�Ω̸���p$�i�)�B�i$��haFr�>'C�Q��>�)@)���U���d�_�g	�!��x�z �U�<�:���B��6��Z�3�s��M�9x".���*��kl�-�۔׌�2�����T��$��˝��U� ��3�M��ϔ"��JQ�p�������8?�{`G�����D�ɂ��˘���>��� ���!Ksŧ��]��;x��<�	.e_��R���X�$Ӥ��c�պ�~Y�ҼC�w��+��� �_˯<��:�( �k.)��G���k�N��}�(l���\��U���ɐ�Yl�����q`�����Wz���$� ;M�?B�4�&=������L�!���Ω��N�Qu���N����Q�/�"�!L�F��H;�a�@_����2�E�+y	K�|bylo$��9�x/�R��>��0*o�e/}}��\�o���+�6[Be5��O�����y@�U��ֿ��m���wa�e{�&�{����IRp6��R!e�vlΔ�{2�����XK_!�1��#�����1�����9VkO����(�n�����EW��5�tŇ,����_�n��*�����{Vϛ�>�;O}���Qߎ`��	~���'-!���Ylo�7w�������9dS���;_���W/�8?l��$��y���q$�F�EJE?ZfM�v{ci��bb�|�ڳLu�V�o�	j������q\L��
�Y�~�S*Ҹ�#�f=>��D�h{�ws�en%F�Ơ3����Ƃ��7��;q!��=�3Б+��$�M
5䠬n~Ee)9s0D򄼣�������q��9��8:���ۀ^l&��
�;���\�DY�AI]��2������N�l&�_��5�����Z�}���<��5��Jx!s�\��g��E~�YA���R���ФG��t=��ڸ��y����8ɴ�(�k�"x��bGZGX��r܏���c���Ԓ���n"���������`������}j^��gW�#F�����H<�C������?؂;ߢ�̎��h�г�K������.[�B��K���J$�ˍx�9f���2!�� x�L(���&鮌�n��ŉ$:F��li7K�ur�-�����',}d*�L&�4Y\ N������(,�<�Se����T����	�@��U��J 4l�mx{l3o���vJ �w&���@�Pt�}Jc�]�8+��1�����k����ۻ�AKu��%��,,�*;<\�|DBL�E�U�@�ڧZ�v|Q�q��;��2;"զ2�w@�P��W�|q�kuiJc�NB�)|�RV�q���FPݷG�;X|V[S�)�t�!p>@�~������n�t�����U�	;�6Vt��׎��Onf�o��T|�+�7�1?��a|�\A_����L�2|LJ"����;#u��B�һԼ^_�B��K4Z�T��g�0����I"������
��Q1#Z/_�#b���7J�Wpw� ����	����?X�)���6@B�e%�>/��ÂU+=���¶(GתwŅ���1Y �����s�l�C��#C�j~������k! ���������S��Zh@�K:a����@�r_NKv��uĞ��U��_?�;���a�i�AP�	�;lș�B$y󱁅�_��cPa?�ԤAFeQ��8��~KdN_����F�v�L��*m�I߳���22�V�T[��;��� q��"yW
0�2j-�3ƪ�_����^�E^�!��;��
���f��Z�>�i̸�\�!���e��M7�=F�'Kچ[�r�0��b�d��^
���4>�3Y!�q[���x<�3�`��F��|���0�a9�
�XO̫����o��s	^�l�y�q&
'�=>1L>����(���M��c�I9_��� i������1�PB�pt���/�i����#haz��`Z�p���5��w=9�bv/��X��6H%��1�����?GR���\�)�F]�-�rx�]�#3Iܔab�V'b4�N�3�JV�J�EJWʬ{�?6c+�Q[8?����N��'\)F��79�8���?�_�F��&�ϧy"]�Y���X wp������k���{�*�Es�)fd6# T��3ͭ#:3+D�`��:��]̐4��[���)�2sdS�d�H�|?<�!�Ո��UM��i��B��A�DyO�P<��`�5!Q�Ʒ���`�
t~��q��-�Vzv*�#��^�I�)|�N�bCp=¾*��T�|#5e 7���P�{A�␺A�b���z|-�ϟ��<v�A+�P�L���ۗ�����K��+B� <�"5���$^�/�1ْs�7��4iW	g�@�ٍ���r�5&�fJ�d!�����1�&�w��PJ
����δ�7�ްq��Y`�?�2UM*�X3��8E�Mc���s:p��A�u�jAROyΉc0�U��t��WHL�o�n����6)<�Q��|�Y�hv���S��թo���݃��B��1�ڊ\�f웃�{;�-�n��'=5\Ԁ�.`�~É8D�;w&��L�0D�tƇ��6�M)k��R���1r�R����x1��dx��m�"4�p0��n��PvYHQ�UT��*���o���V�f�̽_KB�XD��@}��w�PT� ��D?�2��ǩp�q��q G������R��Iq���6�3�:����p�i��ݶ�P�Ա�ֲ~�&���,?j���Z�M���
P1kH���^:��.KL�]�������6J��a��F���#Fx�v�f+��B��$l黎e#����vl���׍�V�;�l�����a>`|�!It���!��s	���_�J�vw}��k_%}ㄟE�鲶�VF���ʽ��~�ޱ~��)Z)�ϙ���O�0�Č���r�>5�75!���u�$�U�{g�%�!�32�	�#�Zʫ�=�e���uh���`Z�˼ӷ�aH�l�	@1-|�&0���o�j����D7̴#��Utx��М�>�P�r_�����O�<�c��-zI���ڸ���kM���-NA{�O��Wƣ�;�f�?{�B�$q<��ӌC�����L��no�g��rC9�c-r;G}�.��_��̈́<��sa?\�ag�a�1c�Z��0��|�#�a�����ff5����i!���UF�i�t�̨��8{��!�vU¦���$Yo���̉����h�R5	��1SL�p,�N.�^ ��S���S��W��s�;�q�pT?�}vKD R�*�-!z�\+���-7h;���g̈́��t�;���Ф@Z�]�$Q���߯� ������'"�Z���ǃRQb<O�����K�q{�'��sk�AU1!st�����1=Вp�DT�dD��+��d'&�X�����$�2��0N%���^>��꤮H\�?5.�*%tm���m�ź�H@���D�s�l)~�:�`��׬r���g�G���[��1u=���2�J8�������آ��Z,��_���ۿ��G*��<�-�Pܰ�I���6����{���P�t���y��k����@�+���_U@�C��,`�	gQ��Sر-�t�l����w��P��ig�#	(!F|'�,ѱ�Ɛ�o_�n�#M<|4X���H��R@���a��T;��39a}��TT�h�x�}:A��0��K��b��gAEcH~5�.���m�m��Ǟ��f�������V$���:9�]a@���z&���� ����"�_:h2�1�ѿas�w���:�wB;}�{؂��}�����ɠ�=DG_�nU���RȠ����]��;���4�43�+	>m� rrj�]f�X�w(�-�/kh&��|��DrҷxE��xϯ����b;
�����nۘ�`$��ك�_�S�0ٚv���;�n�}t֪�PEw���z���s�*s��2E���הr��[���$�l���?������t]�/���8���b�X������c��ˑ���hd~��\ɾ5ѝ���q��:Ax�m	������5K�(�6�K�ʧ���1��L�I�9QJ��^w���l{�Tk=I� ��j>�#��k��W%���U���4H#O?~��<"�F;������8;�,��-��:�R	�m}L%(�>�mFa͂��Ge(s�����dw���U�e�C���jg!l� �� �¡'�/-RK����f�g�\X�'���5�Y��h-���������S9�.o���p�O�)>YNt�g�WYN��2�F~�@�H��:�Z��G�� �����T/�K-ws�y��an6O�l�m^Ck;�1:q���;�| Ps��r�RI��J�ܔ��/X$�+wQ�i�dF�wʀ=燌(8\���:+`� @Ө♭"�\��4�h�/EW�OI&)&�r��7w=��gR!�D�xݥ��$����<~Ź�=���O��������:����4�^Ԁ2ѳ�����F^��gz1Ly��I{Җn'9ޱ���fP��j�a~��6��v�@��j�w�y�_I&���K�	�����" �>��-ʐp��%����ݖ�7Ne|�����'iݗ�\�@ZC��;�FH͑�|n�UVK|�˥~�
�7�-�q�f�z5��A����+���h�N��^C�y�b�0���eFi~|���䡗����y�Q�P�GD�A��@20ߙ�Y%�����X�iw,����z�V��� ?��b"��(��<s���&)�S�J-��ai�6�)h�bC�b�QP��jr��Z[N�\�Y
Vh[ʇY�w�K6�t4p`X|0�u��%163$�7q���PAa1�nofe���R��arf�զW��9a�j|O��Ȉ5�YD��c'S�@���g�����:���Ƹl��P.��������{O+� �Z���f
U�س���תQ�k�ŷ��:��!���I�ۤOY���i���5�R�Y0��P֭��8*{9���t�����-N܆D�t�Tk����� d5s)� ��[�*yR~
o @ǐ���oE��L^�j1Z�2���P�b�XO[�%F�