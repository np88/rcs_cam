XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����N��#�X$���{�^��(iRj���Q��i���f<�>��!悡���yWԣ2�j'�]�>�6�ʆ�[�J�	���B�H�K#{M
8p��z����%ۦ�JvA��t�wH� �H�����7��=2c�(�N������H��u|`�6m�I޷��g��'���Ї�d<`����Rg���R�k

Um����U]z�($�E��@�D�Y�
����*�ͥ��_^ge)��'�r�@^r��u{�<J�g���ce�����Ew�*+���27���'���*6%��Ow���>g�bt����ج�R��n[(&�?+wmi�`�U���4��;ݥ^y ��E������EjD����=���5������Qk^}���K����́f:G`P��p.�s˺
����%��L�-���)T�ib?�1�_��fQ��j� ,_.�{�Y+��t�b�	|V$^2f�"�+~�yCֳ=�L�@���bG� KԟP���oFG��'�R(��hN{�t0EK��kk�#͸��[O�iN�\8{*�܉��rH��0yc��5��en'շNu�����>�)
�-��K���[#9�����UGu6�i_vy�=A�S��F:-=��)�n����������b��|���e��<;�宀-�8PY��c4p�Պ����ؤ�� p�Jv���2�y�B?�K��5�t�L��y�MǤ��>]�,�$�j���XlxVHYEB    32e2     b70�a̪=�>~�L�z�G�t���@^���X�����_:�,;���x�[(1�7j�%@����a,�Bu�
?8(Um��h���a��p�J��?�5��$􌥞�i���l`m�64��?���	ۆA�H9�����ɧ"n.���s���ws<�LHu��6��[�b�>���L��Va?��_W�k:͡}B]�\��އE2m��U���?vX~�SӅ�>�%��8u��MAa�Ox���7=����^ej�$&Rp�J�m��2���r%,S��`�h�Y|��l���u�$� �ߕ���S�:�V!N������
3D�8w�R�[��4�-_�v���>����h@~f2���f������V��	�z	_��yȴ�*a���F���o�N*�4}�6�3ٯ6�nsA��=JtC2dASO�0��p��=�͌�i��a���Җ�]��U�]~!�Ȣ�.rde����A_j4�8��[e`J>�����s	�v�!2̗z��,J�:��.?��3K��[�pO�d�Z�.3�����	�zhv�x�I�u߻��-yY>��܍��
W%mQ�*h���wh�id��U��0�aU0�l�K�NYd��,c2��s�L������k�"���'4Q�g���C>I�sy������Are)�������½�^D��{���q�}螑�Z��/��fl�J�I#	�7t��'*M�wO���wGe��#��]W9��Gm79��Q�.BR��9��[헳�*�#DtRH��Kj}z�&w�iH�c�)���x2A�`o���	�Џ�?�	��0����:�8�1�����DJʿɒ�8�7�Q��Kl�E$�1��FO���\<.l*�e�Qdo���B1�-����$h��V��1Yk��!
�ծ������B�|� &�E8�V�I�,M��
bwp�7a ���ƃ�F���e"��-��U1�E�=��Q�,�i��f�pϧ=�ڦ螇��@7@�����\0 ��7�|�nv~.ƿ^�Y.<�Y���aWe:�p36R�9�c�0χN`c�!�/[@v�:��t�� [Ȥ��1�^��.��9#�ܝ�<ká^5�n�8�:Kh�ܴ���L{��Ҡ
� !A��n��^Y*��X��Y�->)�
�Ia
I��"���[r��=R��U���y�b��7|�cN'��;қA��ߦ���O;~煯D� u�S��s�̋MNUB"���������V��~gC���3ԭ6���f-r�8�s�_�=��A��@o��p��C� CN�U����g��E��J5����Vy����<�>X��NW����ߋ�1XT^`�R���4�t�k�_�9�p��'� q��m5�m�����er�x0b�-ic:ɏ�(Hӱ��v�$v�˵��s��h�u��❋���M#'��p(�l@��&8ɟS٫��B��M���qγf-$9L��K��t%+�k�C�cW>Z��(u��;G�2I~<��ZPL�KS�׉������/�	�C��|��e%��!��Sag�d����#�q7�)�z�H5��޿�)���CN��^__�k��<֬��,W��a�u`L�E��]�gߖ� ���5����2�(�V����\l^o�3.;��+�4���b$����3F����t?��X�>����BR�{� ">�X���r5
P���偾�-�,��n���9�C��1�Xg:j#�K�d�X��.0I��c�S7�A�����ڪ�Q�����Dwc���>�#��G/��Zv"d 2�j��Mb�K[�m)PN�;�����  �QkѡP��>��tGM]�У����&CMa��H7�P� �Ep	�ӪX	�13��]r�?)�{Zݺ��ra�6$sTE.H��٘�~{FR��`�,xI{�b$�2����^ͷ�Я��%H��m�����07�'�����0���u��#����,����kMD;#�W"��8Û���Ued
)�.�~3=]�V�:����ve]Sq�D�����Z�e�A?{ch�^��?�	������$�8�}Ffh����}_�&E�;�Ȑ3��U�����r�B��e��d�g+D�?��c�����˔�qUG>̒�J�=	��������)�3L�.���^���.|5M�W�f�E�%���߶C�6�%gخS������6�J�FJ�uPQ�2ex�IY1��~idlӴ�;�A���j�O�Ӓ/ ��y��⇅r��0�fK?�ݍ�4(,�$ArpW�DF�Gm�9hX��U��L�?�,/���2M�I|��9�)�6�k[L��*��FW�yվ=��+M�EF���~~��+b=�����d�!�G��DO}�)ux�?Q'��ڬk��\�" m�52N��f��N	���AIz����	�Fi����p�}��X�%�e>�?�;�	��Z��Q=z���a%������&�7�|�Jvw�Kq��L��L�{e
��媣�3���y��8b���Z6�[VgO���M��"2�G�*����8c�jZ�y�o̶݉��]� �~-����lӪϑ[Iq�>��gm�����,���������/�p� ��og"�i���`K�ۗ�#�~"��i�0~�5��e �ꀟ;o�iif�9vqEvpWPo�՛�H� �>��7o�
�ƚMݠ�+��V��}fv
x�Y�S�ԝ]�I@ Wgd�9y�5���%sw���%��}z9��*�kN*#d?��������f�y��*_�$g:Ӝ�;����d���t{��|����$�P� I�����:���H�=�|˿�˱nB�5�'9l`��@�D��~`�I��͹����Q$������F폞��m�/Q�9��is��ɆM���F�ȇKn܂kP��P$�ZQɬֶ�V�