XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��k�r�׍3�H9'�Kև�n�Ze��o�
N��M�&Ɋ���}��~^�� .�4"�&�b/�D����xB�b�V@U��6d��#"҉�88�%��P��)���à��=�yA3��UΩ��~��r~�݈
~]��ӫr[�l�>w���:85~r0K<����ʊ����a���_�������p
��a�r!Mg�xP�7��|�^�Kv-���;�|��lB��X�%���Q�(0��A����|]����>0B��E������$��� j��&#�8�<��FCPt��N����p��F����(J�n�ЧS����.�(Z!������<�1��C�'�"�e<	��?(�e��rqu��TdM-�>ٗ��y��Ԟc�ôrz
��e|`�"��i��h�e�<�Ph�_h�j��l�H8������VNY��&����@,AT5�������I�̣���@�LX?��}�O��1�9T]ΠH�r�q���kG�q��t� ��{�m���V7��>[��GH��)������&����o'8�LUS�uY��0�}4�%�g���HHϡO-_'�^����Ư>r�w��*��f�Z�Le�cWv��pc�W_�X�豙S5�W#GN{�Xb�vZ�o{����:����e�^2��r�{��|�'�{�b�ZcT�Q0�4}9� `O7~D�����YoԿ��yM�P���⪨Z��E���_���*�U�˄C�a$Cj3&���Z�i�UÞ���ac�q��[��%XlxVHYEB    302e     c70i@s�� ?�1����㊧D`]G�R��53+$[��E�0��=�C�U���?�$�0�Lf�FS���꺑�QHP2X�f$e�3��i���/�T��Pp洧з�1����!���l�E�w��/�vAu�G�;F�4_�@թ���?�r�s�U�+�0؏"�����H�2p�I>���=���Mw�/�h���[4�ߩ��V�;�[�|Qd� A�[b�\,/}����}vPS*w��qE|���[wus���ފ����)qr�Ն��� �x�*�q$ʛ���t9�k�B1!'߰Z/�%���]a|CX$�Ȥr)���~{�:�8s��pUٌ7a; !��J&���C@�u�4-��m��QnP��V3��FL���e�R��9F�7�Q�Q�\+�n���B���*	��5#Au�x:���1��I�	3��5t�J])$>�ǁд�F�f��[^��d�'��o�b�/����k�h�5��r��-��U20^���YW���W � �������Q Z1�	��3�'���{�X���sY��?Þ���Qw��+p�ʁ�['> f����\	 B!+K�׽�,
t����%�IY��n���� �5�]��� +����"��?����K�7�8ɗwa�&��p����*\볡)��wؖ���˲nE�tͼG��kI΋�e��KޑJdx ,'k�Y�jr�!�����rhwE�=����`�R	�;��,��+�W���4D:���m��e��|/]��/���x���F3o99�[�	R�e�M�2BQ$�)�xk��v�]ANQ!a3�;F,���J̀�>��[�k�/���9����z�N���,E�K�3x�k��SO!�^A�k��BG��[�ڽ ά5��?u�K��Cg!W�j�@�Ȥ�-�F�4�4)�8�Ҳʑz��x��G�svcWm$ ���!ɞK!B����.7�]:��1O�B�0>o˒R�i�{�bj.QY�z�^�{>��������i+��3A�u���kD-@L_�0A\��°�����h�-,/	�H�M�7�ݨ�}ȃ��WC���J^����1�����Op���l��R��c��!Jq���X�V�sJ~_T�f��J\�Ls�"��Ɛ�WW��>����)s�&���.�g����_��Z�A?��B0	�;��`�x�^���ߝ�"�,�~V�8/�u�[6��Ĉ�<�<+;C$�5�z^�L��FHE�yIo�scx������/�H݄�b��@�lx �k`o��!Jk���p0�e����z�����iR_pr��Җ툧�R��H��0�12������q��N������j@^��2�����R/G��E"�s�F������; JV�W��`��ɷ���e��b5:��H��� �-PG�%J� ���@_�� �[존����)ڇ�*ރ
�7U��1�V���Y�(wb�ס^�$���p{����Ӎ|W�	t��9Y�Ĩ�&�3���0�|��ZGh�	]�+��P~��N�bhw�Q��'.��}�q���i��,%�HI0��^��L���B
dw�m9p�{-V�~!�W]��X��ฤG�����c��9o���:<b��Q��.�^1>�s~%]��
�B([�o��x���V�����ї������&m�����.T��+�U�S��  3cy!h�-&���g�Y�1�0��9�p{*k�}�UoѺ�)֐�3�����B g5W��$0[���$"�P\��ĉ��8�o�T�`��ߔ�uO�:a��T�z�n������P����p�hu&�[7t���4wn��G��X�F�煜�v/�,�,���b�`���J����6�嵽�C;B�)D�<�`�Y>�D[P��������B����.�÷��Q�*d���P��.�̭�IH�Ə��I�l����ի=ef��D�7��I��I!f�Cc���L��5��>�f��"��I/�r�`�2�_`��F�;���%��Oc�UN�˷�FQ9���Z~C��w��IW�$=g�@��(ب��a���N^��|�{LJՆ�_��V�Oi����T��A����R�,����l��2D ���ܘ`�[�SH���3�TJ��F�B�{�9��W&�p��@,�-Ig���}�h�)��w��14*�h�3�(�\�#x'�O�279A���\r����%ԥ�p4���/�Y� Es��|�ZUH?m�����<��t��0o:[p�@H���}�����w� t��z�9����G׉B<�<�`g����z�du�!Hq<l�ˋ�?��_W���z("��W�S+*��`�jo�:�q儘(H��9Ur�"�bA�TR��rTﳉ۩�#�ֲ��>$R����W��_�Q�ƪ�#��im�2d'���X' `c�E
����i��KQm@M�%�o~�:��0b�`���̤g�51^]�m�*gK��&A�E���M���uv�Z�ӡk�P����̰���O��ٽ
)��9)ۯ���]����t�i�e�X����[��GD<]�qUb�K���V>�(�AUԙl��D+R���{����fl+�'��(�Oe���{�<�q=�� a���R��a�C�"��p�SH;�o�~��d�
��3��ծ70���.�$�h؍y2 �=���c�R�'��Q��Vѿ�Hn=��Vl�KK������&F�Si�rm2�(�\y4��o���>�KN����IR�����b>��B9��2K��?�_E�Q1��e<�o�!<��-����"��n=F�����^k����>A��9͹A�`��߬-�'��i�lɬv��Z�/�wq��'	�Ⲝx1�[�!�����:�	�LbN��׋���]���3����f�;h���A��J�aPaQ���=�]_������0����DMG9Q>u���[�c|eOA̰C������[hݟ�L�%����V�1���X^��~����+�-q�-���y�����j�c2[�Ț}4�SC�Ĳ:D5q=?#YE�!�F�om*1�B|���A�r�=q�����.+���/�����X���@�Jȟ����(�4��[