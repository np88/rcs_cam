XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���7�W=�@���&�ny�ՏS��G�e4AH��K�@y�\��>&v�Z7�$�D�j}�Y�Bk�\Iz���H#������	V�6�=�p�4����j'��Y��Y���+=#�4�����L�Cu�\)+T��+���1���$`�{�Zi��&��}Lɐ��kl@�^���Qٯ�I�&D�'kR�Ǣ�E���3X���$t��+��A����S�'j%F�,\�GՕ��}��bbA�$����%�oWR���ل#������P�s�q�*c���nr�<|T*�;t��Š��d	3'<l�_����#�e`fIZ6�/�����E�o|Z��G�6�󶌬���s��h{�/M�黈j�杵Q��}HՌ������r2?:ɹ�q�U��k��5��V ]~vsu ��@Ŧ�G����\K���"����Y[k�:N/��_l�肶�H�v�t�l��F��EyH�D�3�ԑT�
�͉$�X�1X�Z*N����V�o�2���M�%7�Oa%���u$IbGӐ!ئ���~J�<?ێ����w>q�d��B��J�m'��n2�-Ρ�l"=T�����&C��U�WTf�*�����}+��ݹ��9h�D!lj$�~uonH���R�#Dɟq��/ ��D��v�.鳈��u�ٷ����sȴ�'fj��6�{�V!%�y�#v�P�\��^��I�K<���2�#]�ݡ��	y���}��zdvb��Ბ��<I[�fw��U��\� ��XlxVHYEB    2df6     af0 �<�0tt�F�))ߠ��n��k	$�VNe,�b@�;Hgg�A�uTk~Bz�Ԟ�isz)~<�&>�m�4�B��f����[��6"�v��'�c��+�xe���#�L�<���Nf���ɡS�&&La����3^��+�����~9��nW�L=��m��
94&�v��3��A*�]\SI�;Sꉉ��ԍ �v�}a+�!8��$D�I����!(9B"��p��9�q� c�c�����q��I��R�j��@��j�
�^;��ċ��li\�!��<�<5H�Z�9o�J��Jա�$/`A��P���n��W2ħ��Y��
�?�����W��2���]~�BM��s����um%i�ܕu��?�Y�V�S&�+�Q%�e"��N2���#��ju����V���Y~'o��ˏU0X�-��n7����(,���LI��Tl�v�p�����[�����Y)�����ˍ<���J�Q��FP%ě�~;�DQ�n�I/"r���l� ~҅���;��0�!�s��8K��4�G��_ZyY�i�{	#���	'HHq��Ұ�����S�� �����ɔ�t��"i��1a���d�;za��3e츞��A���a?H�����rA��|N�1��J{H.�A�D�p��酅��}�v�̉Wg��	ݧČs���vI�A���O_:�۲���~��]1���,j�;١�Ok�"����F�l[9�[^GEfYI��=�ޑ�
]+��k��Q4�<rY�q�<�����{�pŜ�`��:;;��kt��JY*�G�_ 6�4%�%�O��Ӟt77�Q82)�XW��o� �<8/n���NR��*���4(R��#�����~m�Xu �s�u���Q�D|k�.^?�(⠬v��mN׃�A�-�Ċ�3<'UæZ�S���BK�4s}���>g5p���p�>	�%��8L��>e��XT�J6��t'87Od��ؓ�>M�����+3�q*��c�Θ��R��ʎ9�i�j���ba�Ht$���4i9Hw"��M0H�]�͚1�(��Hp������K](���0�΃.�|7���5��q�4�b7�3��h�#ZS�S �훜�	����H��!^F��W(R;A�|s�:QM����Rtw�ڹ���Ęi7�y���a�6�M��5�"�m�1�f>ƘbIt��<.�������<�z8�Ҫ/RI��ؤ>��>�_�����p����WO��s"�-�
�����c���#�Z.�8O����/_���1��).��`�.�,���E;�_%�\o�#��)�v�Ӳ�j��6#(òC��Avu��}�ךc��Ȼ���L�|�NW�G��C7� �2M�co]35��=��]6�8mHc����Xrd�-�g��r5��M��_���ƥm|[�g7�=jG��bB?�;���~zTYZ�>��t({C����!`"RO���Z��"�=5.�y���!������aM�wÓ�(q#/����DH�Y��N�7iK�QL��3�҅����H�}h�_H�C���� ��{A�k��4����Ih��!�X�L�Z^+��0ꇐ�J�f��"�"�w-����+n�_1Zx�v�J�&�4�UzZG�;���#�9ȋ1nH,�pqw!u�C0
*�/c]�=���T1���O��e��SGV��t)\f��vg�g�l��pJ�8����M�o�HtO��m!8d3�K�81ϜP;�]1��J��'<�Р^z������d���pj�-H+S=	�̡���b����F�ȰP��j�JP4�h��/��Ť-�ec-&q��GF��F� \J�d�*�dC�BU?Lw?�a�x�JROa޶���C�!Pɶ{�_�x��~/�X$�D����{��(��(��#�~g��Dm䑈8N��T����P�9��/�^�u�2k,�)�)�.��g�b��ZϝI��� p����c���捄�k�?��Z�B��q�i�����g.,�2$�B������5�<�(��0T5$&�^a�F�8g?�R]���^�}q��Vr�f����g$%�����~{�3-��8/ zKeg�"�67�.\�F�����l���*��7���"�y��9gg��c��}t�w8�`��m'oW�h�?`��9Ni��	@c,�-�h'�
B��G��s@IR�ޘ��Q����$`�LՈm��� �����<+eI�3�*�0ß�����?]E�Z�4#�7�>){�Ɂ<V��^�C!lK���%�x?��^p��bh���$Қ�P���7�\��=��[I�/��3��.��rɴ
@��~|�����0l�H�t8�����2��4_�a��)5c{D�4��A���@�� �� ��ߧN��g�c��7�YG�G�JOe��p.{Z����ѥ�I��`Wn��O?����#Wx@���G����3@����+�أ�%��7����d���&��3Er���uĕU�&&�T!�靖1�����1)N��Ia7�q�Ŋ4v�T�n��ǱQ{�^��y���ߞ�X'<��4�����_��4��>�s]0'�zg�7}}B�4O(*\�l(����U���k�s�g�K6>,+�,W
N?֙iP�i�s��,� ��xh,���u"��S��\
r~���ڮ��;���\�����3�f��ъ�<θm(�dB���7�,b<0�?}�����H}��괅�O�=�[�������7:5���
ڲ�� ��jy��e��?2I�� 'v,��gլt!