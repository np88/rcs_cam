XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���q>�"���/\�xOj�@�-5��9�ƵD���\B	(!,�z�d%������xw�Z�j2��1A��>u�~�m�<����C\�#��Q����ܛ�@���*�(Pܺ{Ԯ�B+�72��,1�v�.[u0�/��Mea��x�*��u'��S�.���<�(9N�G�3�<��溺����Z�KXxi^�C�I5uu������y0,E�����7LC�<�
r�J��+��%.��@]�����M{"j³�V��H^�`z�v������iZ�&�Z�~�e�D�|�tʻi�y<��BC��(���)�}[�X�d칎 ��0�]"��Z�z!��au��˘�Q-�Iܦ��l�I`��'�.
 �� :�zx�ϴ�%f.�_K��$a����O���#���z̒���UԷ���F�XY+g���)���#�B+���)��&�ln� 	�1�,�f�?o���� �Qu3(�*���n3�k�]���o�¹��1+�=±ՠg�}0���*������LtU��IM��B�&'�#�x�*�G��B�f5��X�mz�x��[oq�@����nwDzY�Cs����2t����E���6��dv��J� ۦy�M���t]����(�<�
:F�t~�1"|�:��D�G9�yj����d����̭p|q��SSy�{�MI3j@�R����Eh{�T� _=U}��k�j�J��\$�tD�Z�<���R�V�&ޜ'��r;qӰ��%*��q����ՋXlxVHYEB    5073    1100�.�"�(W��8F�C�����S=�Yڿ�&Ǿ��ˌ���t��tѓ�j�s�� �VS�~�'PG����+���Z�\���pד���xR��?Y{;�s�%�
�0]@&�՜�wm�I�_��]�<��;�%^��	c?z|Sv�|�J�b�/��n/ѓW�=�_p�]���Da~����~�ܘ��!Nj������!��M%+c.�9���nQ���Yv]V�E��ߩy����-�r�=�f���yww{�}���-0|������e2���0 ��P5f�|6οG���lXr�`���k����z;�[>���<���B��*�z���#.|��ױ���U<?�I� ˀ�{�LM��F�6VHi�j?�M���ds)�.��b�ɫUމ�J�=�qƱ.e��	���tb.��3,�i���;����K�$D�?�rx�U�0wU*/�X�B���T����N^_,W|A��փvV���U>J+�aY�� ��҅=���$=�ͼ�.	�٣�����W�z�R�o8�F�j�<zCW���?_�"~�Z�疹����z�Vi�2�2� ����N����6{����i�����#Fb�!H�M�r=����z�����O��Є�񸠷�Ob��Ԡ���$�JU�c��P���S�$��	�i��|֤	�/�aa>���k_+�8Ͷ��)	�`~Ia�B���bF��x�j=�C�A8D �	g�H��T�y���[_/)=.��	��nk8I������V�� �����	~������J�a�������#fұM��[���ˈ�=F��+ �#�Т/�屭�Wi�Y�z4����@�&6�k �vW���G�G�����=��]B�&6w��D���r.
������mb��(�!�?�r��P�WI���㎭��`��{T����'j\�	׸���nx��Q{.5���YsW�I�V,Z�b>��%�F��U�sS��������_F
:�GEl��[�{�ۙ���������~q���_�#�j8?�O�N�d"�<`ם&�@L^�K�ffK�8�ԗ�F|xAӂ��?��0�3x3Ї .I�wk���7�g�rZ6�����;^�&�W�8�����-�O1�{�\��?��2	��5�h�-e���Jwi�:��5��"�O'6��t�l��Hd�u������{U:�F�;lm��h�"��r��Ӑ&��Bc���x�c[�����/6�C7�p������Mg�̈́��nA����f�+��J<8{=������E*�Ń��+��ʯ��ޢ	R:W;����'��9�V�I3�j�-���4��4�ax��n�/zi�l3 N��J�/L���16�eH���'���� �!��$�/J�������j��#`���!42��w��]��Jv[��'޳���0�t�P�Yz��,#�)z��S��(9Ls|OV!������Z�lLnɸ�^;jp�D�j����PB�s���kE]�yVA�,���Rr^�32�O�֑P�L�AW��PԔ=s��/����XXQ��~�Np�:����,Zǋ�fTW0��}:;�v,ti��#F���V�6��ge���.zIe;������-O}���Qɥ2V1:V؃��+��.K"���{e�_�v�2��Z�,N�p�j�$�<�6vw�� �K�����U��<P���P�r�eM��t�������~خ"�|�%��q��n���<6@7;��j���X�^4,�U��/���a"-@�)Wc���{7X��Zwq�����+�jF������Ousqg��8�낼,W.��)8b���3#����]��)�ۭ���CB�)n�0�!b�Q�sfAn��0��x���0��CY1�U<Up�}�I�,['ǠⰜN&�����f}�C��2������<���SM�0�l�X�[@�����t���P4I;�-�34_G$�-�BO�2M��ٗ`Ӫ�Awe{3=?���Hy.u�ok]�r�����E�n�W&�?������u�������g��G�i7�R�3�b�-#��YP�,t���Qq�i���d��{�vv�*#S�=FW)q�V�EW/y����
�]��X�.���ӧ�"nF��d��q�@��2���y�6�8E8��[_ݗ�3�����pm�����;���w:ϐa���5���E��d�DW�i	/��Px�;�Nm���6jU ��H5��޺�1�9�(�>�}�+�G}��L��C"W�闄����[�WI���Q^49bq�Асg�͜�[�,��fb��~� mΦ��=*eM�7��D^��	s㩄��B�ݟ1)���	:���.�=��۟���t`�7�j%B��A����b��`�61�6�Ŝ��"䩰0�T���J�}��l�L�j�~�h ���5�a
Ț��.P���\��S!����E�0t���*�|�y8uR,�L��XuE)�����C߼��h���57���J]L�w܊܋v���n��7k��	���T�́:A9���/�2�P��m��`�/T��*:5�/?�5�~#�j�g<c������u瀦]?;6v�V���l�g(�����#�.�E�B�ach�H���W(P����$y��z� �̽¹OD��f���^v��{��"@������z/�X@l���ji��	L?�� Ze�O�!l:�7F�6hn.O=�ꑦNj�6iM�ځ���j�`O��8�C��իC��t�Q�N67ʓ{��fZ����Q)��󟿛V �|���0�1�*0�U��X`�xF�D��PLܖ">�t]��b��!�ѷ�:8*�I���o�P�K����Gu&Z�Iq�q��C0t&�#4�\���2��������Ut8��TX�Kg|#}x��{�3O�)��W��QŢ�ʺr��3��Yf��`�h��[80lj����QԠ96TR�e��wB��C`ӽ"����10��-i
��n��=b��4C��@��>��)��Y��N>��E4�&C�|p���������XlȃHX6����d���V���!�:�${T
Mp���
�����^r�̓�j��o_L��^$�ٖ��S�_-�t�T�^"��PM����#�5�w�Q�=̬Ju��r��l+�^��mq�0�"<@��`ѵ����EA�K~W�~68p��,]��5�1�8K�\'�r�$�k�h<
�,�N����Y#��XQ̶�As#8n*S�Y��#��q+��\'7c��%��=m�ޫ�!��y<��nk�S������0�f�3m��9����lH�����Ur6����=W��%���5��x��kj<![*��ЮX���{2k�M�����yQ�������y�X���)��~�|���7=�C3'9��3U1�rI�L�wϏ�YA���nӣ�Ԕ�*R���1�"I��SԻ)��7�x���Q�6Gn��SBɽ�f�M� �T�����J>c}k�v{`䵷��%k�)���ר�z����s�Mdqv��;K�*٫1Y�IzJ�"�;�]��q���&��)s0x�B�c9Vz꽢X��2�Q4k:���V�S��$��"pB�y�xNZgcr~�l⧚X���._g��E���_�o�$�T��D���!����M����М�zO6�3��/��jqD��z*�qN�Z�_�FNL%���PE�m��0C�������t��D4S�~ť`��w�o�oc���4�+�f�Jt"�e!����f�z^EFO_S ��v]�p̇D�$=�%��3gɔr]M�Ђ9�ZX1?��d��^n��§V�w�Ի0���q�5�vŷU8��jb�>V��`>���+(ƂsP&�E#� j���eAG-�,��:�̑��;�-j�пХ���g�b�o;����@���:�'��N%�mX�6k��m9�)'yȿ�p�@"��Ј%~!��Ygp�	������}�Q)A
 yxu���"��֧�5E ��F7�$�V��-"��`����3����nl7=�q�Fl��&E�g��]M��Bs�%�,�ڼ@�U�*3И����*���5qy	y􊽚L�Sm���?𲅣���RT����5�A3�o�1;�2�ڰ~���F���
HY��8��O��烢������\p#�1L�o3T3ݲ��:M?������i�7}��k?����+Q��lX��d!G'qu*}�dw��1Ff�pؐ��AD��8�M�n_�j>L}r:�#���#ujG� ��f!I�=�Z�