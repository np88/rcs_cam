XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��	����2�%�{T�4R#W?��S���`%�5$l9 �;��bk�u;�e���'��X�����
A�k}��(d��f�KIɤP�}+��F};��8���DM��QIp��&���O�o��ܚ���4�P�TyS���{�� �2���\�ش	�����[�3��3bʘ���%��@jMz=*=`{��0H��3-���ƏA�;іJƻb�����L�8���=�k��f���4��Yy���}@���$\|f�Di�u0�|a.]�P��y�Ί~t�Go����g_�N����������;�*n�q��D �Ғ�Țg�
�4Nc�/'J��gk���V�&� ז���@��V˘r}�$��gD�W`�m��g;�y �r\z2d�m�
���(�~�0�Ә�Ax/{U�z�|��������l�.3�ض�Y��?\(j&�!x����Y0��������!S���M��[�q��`�3��a��f|Gҡ�1��I*��(�f^�v��8P��$,ˢ�Nׂ�e7�4�4I�̃�&3]@q������jI��Ad��#q��y�[��F�_�N�Wڬ\$����;C�s�@�n��ϫ]���
CM��@�w�z��.�EX�J�j�*�C�u�i�k�:YT��t�Ä]P���-e��^p��!*������Z�շ��A��<� -x5v�F���Ӊ�t��q�a$�}<�2����W3씒<P{��M�l�N@�xf]��.�j�2��#�XlxVHYEB    aa31    1e40ꚝ������V��l&U+kֳ�j���{7�c�U�袆}JV*e����^-VAI�1�Q�-?���
�N�`S����zk���U5�ʿ�6�D�n=�[��6��7B	5��٤������0ѳ8�yyϯՉ,Đ���>hL�@�e�g/������+T����"��e����n�&����rv�ԙ/���7�b���M��k�@o��C��c��*�~��[�<�B�L�D�5��f���B�#yu��+���w��c�N�O�Z-��ؾ�t;�"v�x�M���C�F�n�Ft*UV0g�3q�(��#�/]C�R#i�׿���n;#�34ƥ{��ȴł<}P�:��P�z,�9>D�"24��T2V�% ����چ�"ɦp�t��� t7I"�F�L��|��"e��݅Y����o��姃�=7��h� 4_a�}k)@2!�
�b�5r����4DiH��]\җ��4vK]m��<�v��P�$�r�q��\+�E���I�R*����.����8C/�Z%�����Z�QrX^����VaE3-$ �R��O�E�R�~ĭ*pML�F��3tt�)gF�[(7���k
y���`Q)k�?AR��Rq����qV��_;9�)�+(rE��?LAa���%����W�˫�G*J�ݚ����Ǯ���2����_��~%Kԏ!��)R����y�����Juj���{�<3�����}ڝ�,�Yb�e�F���?5� �:5������Q�4� ���V"jB�$�G�UG��� �f
Z~A9a�(É�#�A�l��s��"�p��.��A�"���r��a~dm����oWz����D���7s|�|dUY��+���	��u秂hGq��Wٌ?��Zp[��;�>h'�����a嚁�#����`�
>e�k+/��*qxڶ]� �s���}�Ǥ�.�
���A��Sg�$2�(sN[?��^]RfN�$�N;i���Ѧag˜Z� ���������W$��pB�痄�ve�87��l����|$��82�5Rr�\���g䛻#��/Q���CDהWz���	����b+y�/i�-gX��T�H%61�R�`����8*ĩ�3Y�5��;,�쇺]�BO�XU��3��dP���L�"�
r\Y���GV�~de,�J����~����ӯ������G��=�f��Dei���4�|p&�	�UK����*�(9��ڃN迯��-�{c)Q���S�z�X�P��H��,H����	��P�-V�rg���ŕYv�φ�g;BUECƎZ�?�8�zAA����2��f�V�Ϸ��i�����K>\�!9F��	�+�s� �W;תac�4�*?�o;�|x����3�?_+Hr���~�L�����2�����_�1�Y�,���Qs$���J�x;�������t��-_��-�^�V��g��n@O����;C�o
m���<�	z?v��]!�7P"�
��Eͧ�WS9i9XyĶ���zV��V/��{��!_�y�gX�Ǝ1�t`�����<I�fp�w!�W�L��.r�ݍ�4L��k�i���Ok��^C����QSmr8�oq�.0��BS�r��0���pD������7��0~��$3�Dn�9��\N�,�)��~3��Xl� �F�]#�e�H�A�~62�[Cj-��w�|����99Y�tѽ<�n��N��t�3��}0d#�l�r\���'ȁ�J��R�<A���wzm�׌�&P}�uߐ�g܌��r]^�g� &�I��,y���� ��4�Q=�s[�s��#�f������r��G]�/q��Z�.GZo�5��S�E�Ep��H�>�d���fT&9�'4���;K���M�hf ���|X����P©��k	n�h��/�B�~g�+�������P�b<�58��L{��vSVo]svz�U����SÕ���f�H��*�Ϡƹ�=N9����"$���ە��.FnE@�p�z)���2���	�4]f��o�#]+��l��J�SL�����+�5"�W�<9����_���H%�x��dl�^�M���<�	����ix߃�T���;�Q+���X9a%k�;�'��W��}� -�����o%�W�y+sc�=k�5��l�09�q�/7#��.�����?��\�9}iy�U���c�_)�)�.�~�j�P���V�q�D�����1��h�_Z?�����*&�EB+����v��~��!t�f��a";2�9�1�=(,��(��i`�ʷW<��2�
�	��A�q:�S~խ��X�Q�8H2 H��R-�ْ{*�T)g��n�BKY�Am�f�L�x��yH�|L�	oM���5�PTK�^����񢪊m3S?�v�С"�e�L{�.?�"FR稳���v�h�}���}�{&�n���R1R���R��=#��ob-���8ZxE����L��Y�/m(/�X�E�{��Lџ�ø֬�:��?(���ͳ��w�xs�m�6����b�U��a�R} �u�3��P�V�J��x����6��L
�D)�A(pe�݆Z�qDO��XFo$c˼����❒6��[F�x�;D�~�+��,��]y:T��;���O;�$���N����@껔�}�uay9Ҭ#���.D����=Պ�(?I�Pv*���z�������?H��c�H�ή�����E�	���+�k�뜘�P����_���[^��h���8A�M"�Ma=�Gd w�2IW5Qy�������" ��=X��CA0��_}�ĉ�����4<�PN��ZM���C:mE�dVas�x3Є^bg��S����Ba;��k�!8@���h2LX�ɪ��'CyG��� ��s���|�� }d(�s�5�eƉ"��N�F��uȺ�� ���R���s:�<������y���8yT���;gch���i�x���ތ,�B.c��V�
"��2ȱ�L��A����u1eq���;�{/E\mۼ
���{��QYi�* G���&�?  k��5i6s��/r�v2Z;���s��q�;/�f��Mzwƍ���|&��,��Vm�3v�cɶ�?��5�N�-�e��������Y���A�mu"ȜQU<��90 ��F=�A�D���,��N�n�[J�.gZ���[�k��B�"�E�}�e�"F�Mgeɟ��X��}�1^a�R(��P�:/~��a:\L�[&'�j���,y��8���V�����|�& �H�}�0��muK��U}�Û�<�u��7-�o���x�^�#��:ʃ���g�naM��aaƾ�s,'�FE&v8���Zb�0��ߑ��3�Ղm1�o3�Biࡠ�^2���]��GW�o�.94־l;e�	��e�C�][��M������8�����Q�.H��>r��]�(��]r�k+cի��� Ji�^!���F�
�v#���<@���K|o�y�����,_�T�#3�<P��<ʭPEA�@P�J1��ӪI��8�{�ǫu�0��e��mŎ��L��n�t!���B#���Ps3��5�:Cֆ���|��Μ�e�y�C[rI %�s�~�+�ފ��,�}_m��8Z+K~��)�>�}u��,�����i��c�sF�L8e�^���Ļ�h��lv�ġ�;��g���ǑX�#8_�"�9ջ��k�,�fD����w���̡�Oڮt&�\]#�u�@p��>|5I�-�7z=,��t��cZ��Y<��7 �x��(�.]r�ҁm�P���->��ے��Iq��l�ҺP�2��c���	�?���%����/yk��r��)�3�9���V��r/�!L���Y��KF]�ZjRa
�P5/$;��Zi�D��.\�����L�q�aU�*a�Xl���8M�̴�)�y���C����l���f�#�z{�c�z����N?s7�D��\��K{��41�Q��ӆy��t�qˏ�pu�A��/s�G� ��DI�+�4f�#jF� ܹ)qź|^sr�����H&��֌v�.���J���?�:'�4�d�� ����m���#i�ה1 �=ֿ�Π�26��_vǕH\#&�C����|���.����D���y���ΊR)j?���!��Q�:/�(?�%n��ݯ�i������c�D�6u�~i�ܶ�]�:��@��R93�0m�v�o����E@T���[�!s�aZ����
5�؎GSyT��|>\��1J$ﶴ�a]"��d/y)R?L��Ad�(�u9�t<N\M�� G��3�+
<�
=ة��.��� �PE}/3�������4�����y����a{�hcsqwGlTE{����Ē��K��N��sr��߆��?GZ�)�؜���H2��	�ޔf�㄀��>�⁄���*�dl�����5dO���HU0�N�����H~b�A=��7�-Y�����_��G��\c��A&�;_qD�V��������{��Lwi�m�򨊧��p�l��{K�^�ǧ�N�{���tnQ>�GJ�	-M�Q��ʍ������H�o #�0����e�N~�1�=4Rr���2���<qB8u���%
�5t�Gs�Tw�Q�����]5��uCNhj��s�lˀ�ͭ�Ǎ���C!�V���"ڴ�t=���l7@�@һk�&=O#�
�%��cM���ݧ�R���i�6b�h|���?�U���~�"2&�3e#�����.�S#�
W+\�,TV3D�w��R�.�f�ђ|篲�K}X�L9�[���'C(��`�ք�a"y�*��U����v���{���(��F���^��H���[8>�����l�<�5Zn�X��;�N�l���}��ch����y	0��⋣�E* ]@ݻ���;�Y�(�ժ���u���^�J��	ݰ�͏�i0��4C�j���k��Q�_5�0yGe��7�3���c��i\�M-�&��%B�@f��r]�vQ_�ؽ5���3uL�~{_���m:��������]�B�Eǲ���5��2e�ך�lmt��y�q�*�$�[�Wy���(&F�{�K0Ϝ�/)�3��2
�	U�ݶ6�>� Re�a�|/�HFPe��% wT�r� �U�����M+-�RѺ�+��,Pz�	���)�n�2�8�ZѰ%(!�������iڒ\&"9�$,�#�����-?W�r���"jq=���B�HL�`[�x�u�G�  �C�V�M����y�L��FS���?s`3�P�M����ׂRV�b��>�}�?O����[��̇7�Cv�����{���nZ�{�">�a������|�9LZA�U�1�s����O���MZ�ws������'$Y�L�O�"q���n������e�ga����>�����|�$L(�მ�6ljI�]����P�%�i�Y`�gU(����ppzȐ�d�����z�I��d� L7��Xx�(G���j2G�\���U�f�@a��J��N�ܡ�8�����f��CE9�����,��ជLS�2�oR�/�|HЋ g� �.��m\�K�,���mI��&�Ȅ����D�hH�U�VCdET��#Rk;�/�m�Ve�԰Z�7¼�rL#�����Ra�O�8j�b+fäQ������g����d��1\�o�=@��y	���UzFk�;�SB���M����n0r�°����ސ����}۬=�z�6��2-�I-���ax�X����i܇'-Ė��Ws�B�!Η��g~5=N/\�Th9븈��jR(�h��zN��fiQ�+k9a��b� �)Y�i~NqDf��4n�kq^wt����_(B}$B������Q;�d)����ư-����9���.�S��z��Ӓ�bja���p��K�q�; ��k�Tv�^C��Zzb���z����Ja��/����4\���?�BҴw�5b+��&����d�kh9)�g\���SJ(�t�%9�#n@j�``�NxTX�l~-ُ �W���p`1�w��@1Vc�^X���(i?=� �O4��G����m�0S+r��qB�^������vǑ�}����L�Z3A`5�=f2���ZCy!Uy�R���W��^e���Fb����ك�*u0�`t ���w{����D���!NoEJXEi�Ƨ�g�Q�
-+�>���"`��[F�8R�KV�g�aU$?��>���$f����s>ֻ�U��=$��L�����Z�����s���m�Z�6���@n���2˷��@�mA0�D��l�౗�۬�A1;��lݰ�(=M��r��Ed(�Uv�:�&�b"jt+#�����IG#�y�X����sg�W�D6���TM��yl߫d���ռ�7������tp�B��.aSX�	�����r�����g�80ͥ��i���G1D�7~V��p`w��	��]��|���$iG��u���-�J��Y�&!1��fOnP�HG��x��I]#v��E��˗/c�1����.E�?m�R7U�9��-�f�f2����CV�U�BqI<�1@P�2��*"��Ϧ��{��ڧ�I ��}��y�%Js��#�h��A� ��lN���j��#y�<�fF�D��>@_I�A�F�pL������oP�OXH�0T�FZ�z�� �VAR�Eh��� D�?�X�۲���������$E��=�}.�\d��~j/,�%��������>������G
&l*n�������ޒ�W��c�(�)<���ݎ44GH@���fF'n֌�e�Z�������	��a	v诶����� �G�@�b�ӏZ�x��ь��{�I����k}��Ĵ�1��W��G��@���3��ު�~�2�)Z_���W%�5c��\���Kna�~����!��W�vڭ�E��p��+��*���L�`���s�1
��e��ם���Y/;k��&��~��31��"�LF�m��KE�����g��p�9�*	b;C�I` �WS"��w���ˀR<4b�{hgx\�o` ǳca�bs{ j=N��b����T�Q�
�(��A.�QG/�t�-;������レ`�%�"�ç�t��%O�m2o J���$x=�n'��-��%��Hk{b-�w�Ct�֫��o�ݖ�84~U�/l�����n�a�v�3hL�ڿ��^�a��x�v��5y�g��Y��b�qn�,�����`5�$�t���Eq.�OW>5� �I�y�ND������D�H�?|;��u��A�A�z9@�;��bo�2.` ����[M-���@2������?87�2uOb��n'L�R8�jbd��S�R��:
z.J�a��.Y�7.�iԫ��}���V�^ߏ�Y/���t��+t�2�v�pҶ���r�`�3��eߞo�sg߀S�sT sA���sg�v��[�f��N�5¡N��%�ئ��ܳ��buN�\�I2�m����Bpn�35v�\HQ99j
�\s�+� ^�c�gGK)��a9 �h���m�j�jk�����ꐶ��� _�}9��[�*��]��ӑ�w���J�h}�?����?L(b|'
Fo�����v⾾��3"5U�c}�ӧ�sb0�ҫn"t3a#