XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Ɂ\�,a,feZ� _������"݋0���� � �K�;O�X'��=�W%�7��|�Uc���j�#�4���=��"P��*�i�ja�C�)|.Ѱ�%�Y}�:��X�τ�F����A�3<� 7g/�✥{�
� �Ya���!�1h؍,l�ޡ/�*���'���4�D�B��"Q9c	��"�H��f8�#b80#"xE���/q�j�J݌�I�G�xA&-*2�F�&�&T'�Y����'��2J��I`W2�K�!�5�-�է�h����#���60������I2�� q�	Z�j�ײ�Փ:0}�����E�_*W3��G����4�j�Jhw,辒U�
�i$���`����f��H��Ԙ�H`���$87�Y� �3��=L��F�/ ���׸�N�k3��7���^�q��8m�תRW#fg ��D���B2�Q431��UU���b�8@/-W��-vܤ���dɐsC5�v��;�T+���K5�^���EP�l�D�^�.�M��1����7!�� �z���e����LܟZ�խ�y��nԉ�`�q�n�����&����͡X�)a�9��^)JHr½9-y�ҫ	ouXYj{u폒k7>�Ή����-�;��d�~7I��� �mEݢ~"6�� �.
�'w�g,�PG&e���O�ȃ�1#�]&l��a���g��>�&~M��T�6;H��$*Q�[b�ɥ �d���:Oh ��	��dl�&+�i
)�sXlxVHYEB    63ec    17e0����U�j��Rְ`B%����*D,Ju���@'�@������x5v ;�"(�����s��cw.�.�C����J:L}�a�kO9H1&$Uo���u��p���Ujy�d�Q!�͞��5��QEf�mьh=N�*��|A�Q��w!W�*��U��t:��E�4kI@H9���)�Z�A�N��W���s�RQA#2z!	W�����=ʟte��aF��Rō�3����D�wrc�V��ګ���u���}��?�p�� �鏙]yN�p�4��,p�ؖPv*�%��?Mƀ��9y�"����ꔮ�?&Ăo�|�Pј�,}�L�(���r� ~;�><��H�y�^4���}/!Gf\k��7��b�[>��|L\@�-!�e�iJ��$վGL���x,v�[��ԇ|�+ɍT�y���O8�0F�ًb1�8Ӥ��;,��~pɴۆ6��Ȼ��9���j]#S�̒T��3ʷ��=���w�5��	�����0��`uu��z����P��o�!��� �5�o���8�MHR�=�)Y�kt�; �!�ĭ��1C;_C���Ag.�.G
`�P��,��C0����Å	N��d�-��Pd�O�+�m'7M2�q\�`�҅�e=X�{�"�w��9�n9�^�+O�2��&=�h��b~�y55m���K�@a]��?�	���+K+D4}R7�`�/�5}^�-L	ͨ�?L����:�8��=<9f=����RL�q����0\��{OZ,�O͂ꇮ��4�~�,7�^��fc�Z҈z�=G��jP4���}luF�Z�D+d0	�~A͜���c,�1���}C����5���RVv2���ܗ҅��NX��R�Y[#&���c�&=��l�lC!V��|��d]�/�!��S]Z�%Fx}��`�a�5ӗl"���:���-OH�N��qF�� �wRx��K��-x'�)��&1�ާ,��4|�Z��I��MD��)񨝁N�t%1�З�Uʳ.
[���Q��2���8r�6������x~p#8��/�Aiz���6����|�y�OuD}d#6JP�^^C1����������!\��ԙ$1��j�DA��J���\K��xm����}=�t+k�H����d� ��I�k0[wcg5u�iU��Y�U�ߩ�g���KI��)���֩�X�`�~���gϿ5�2cs�C쐅�֬f��г ΢���ն]�%��	aaS񃇫e	h����Y���������u�6���!񦈲̗�բa�u:9q������%f�{�I2n��#�����h�e�r�>j�<�L4`06� in��i2	s�LQj�m�B��Sӎ�!�:z-�e��� �ϔ��ܰ�r�.공/)�G7�� �RY� �$�*�0���b��ƙo�����N�MZ�(�����"��p �(��C��˼,.R�#M��O�Cހ��O��������;r�MW��l���`��yL�l����ıMb�/ʈG�;�?���<ߜn���4�T��JPh<��`��I�U
݅hH���*�@hh[E��y�-�yRgZux25ˊ.�� ���&��o�_(T�h���75Z҂�4=ܤ��OM/.�~��,ku紦s���H�
�]��:��=!��b��,)���$ D�z�$�ka	��i�E�������\��̥T'� �d:�75sM�F�%�B��Yҫ��m��tY|�
�t�`"���F�]��y�����\�G���h��e+���:b��c�xo7�������ޓd�yW�N&��D.a���y/�N��s���<T�<����ey���.�R��p�$D�-�b����g�l��:�,]Ȗ��Mv�b���}���נ7.�v�nG�P��_s˹[Ć�d�թp���ze�L(H�ؾ�<�����p0��C��q�9�����⶝ݐ���м��e��Z�����vm��Vf�a��s�Ò��B�|�~�k��/��V�3yل��v�L�u\�Y'�����#2y�0�b�p��g��	M�G�M���Bls"$�O��]�uӔ+���; m���:�A�f�����(�@�B�Y�q����l�fŻ#]h�}Ї��J�A�r/���g-�����
�8�V��Ѧ�LA�9umIe��r�P�𶱟��,�����j��"4��J����"u�>����m�IY�����h|!�SS2�`��p��c�}65�7:Ga���x�$��+J���a��d:e]`���y����\RP7�c�s�� X�M$9�I�s����H�+Q��v�6�����$KÊX�&!�K ���7��/l�vwv���g�>%[�(�j�����$[�e�5�c jFY8��<�t���Z: 	rA��:��l��Ns��At�����x��3��Tl�L/�(���j�4k<�6o ��1�݃�y#�\9��=�O&��ì,�@~����c�XLo��v��P�?l�����~�#������M�D�`�}�.��D�gm�&|Xa;�(��	=�������	1�v�����Fq��gk#>,����Ga���ݿ,SXr"
0:ė��|R�}9��Z��dC=13lg�����`��Q�]�Gw��d�{a 5��/õ�a��hfz��~"H�÷��QJ���e�@/�/R.w���IL}
) �:M���&�8�?Z@i"��;o�pd�7#?*+ /�C1�0�ɦ���YJ����vR��"sH[HzΥXE�M���g��_���@��_�e�v��%A^�����lGcH;9��nW�d��!o�ʀ��w��
�]N�5<ht���E{�Q�z��P_:)>}���'��W����{��8��m���չ���H�]�ږ�����Z{xՀ�� J� ���.�IU(��>P�L��DG��A�"g �>="���Z�ΪU��Zvs��E�F��;8��Q'�{4���GL�n�(���B��2�f��������q&
V^�(c���4���q�0o����m#���ƨ�����%�]msO�m� ^v���F��B��v����A�L��?"�����p�;$m���Ie�Z���x��`�޻w�h����q�T;�������K*�M����;+�Z����ۭ0t%�ڂ�I�ڜ�>���5bx������O���Y��������σ���u�-��27��A� ��-�%#i��9�X���X�e2X����e�i_toX�C�dL�'�[������p�/��K�B�]F^^�5m�1jo���,�oh���|�Ti8fß��H�(���A5�� pWɕ�䈉h�Q���z֢�J��ͤg�Ѝ�B}r��CM	u������j��G�焿72�I������Ac�Ĺ�|��L��D�����p΅z.M�@D�9�*B�A����+uŌ!U\�����)8�����1f"bm��3'wW�92��få�-�ҁ��.�^�{GV���P��H��c�{�L�����ɧ6�y�^�QZD�eo��N�pZrzqy���TU��)m��;�ILn��������K�?�1*/GaN��¼ËH�8���v�����o=٣�ٞ�N	��,ğ�b�� �Jd�����G�dF.a͗�ԗ"���0�ܜ����ݚ�޲�R�=�U>�G�"̂���TZ-/���R�p�E@��*�ك��u��8ܽj�U�t�_�յ��O|#��&X��0�+˯�.D]�A1�Kd�	 xR)L��}UXT �3��ed��Jr�a�y�zO����Q�Z>]��`�5zd|���F��2�8r���&O�D����`��M.���n��4e�}���ob�Դ�h����b�*Ah�#��j͌*�>�;���=��
��HH�̼tn,�,l�hl:T�G�C"�B�a8;�<5R�<���TF�L?1�� \zc[ݱ��V���)D��@lS���
�ŉOق����ƪ-+0�2�.]�|��|��4�[�+��U@}��ݯW�Ɂ۲�ϥ5���}�=��`�ˡ��̓AV�)���e�����D'}��!��z�嬤h���mn�H�
��Z�і[x�O��=9��~�:��'����wH&[ ���'�Id�}�� �)NYK�
?vwܮ<�maXmE�,�"�,�q�v���O�3R�[]�&���`yS��"Zڰ�=��Z�y�7M�6hH$�`��U1�:���l6�����>?V��J&H<���&�s�$��8+���9�]�4ה��;�NС��Hu�j������4�׉?1(٪C�N�0��ko'S�.p���[}Z�QK��������
F��aE����0���Ј��;T�˄��%�v���8��_�瓷CZ�;�pnDh(V�����u��V�e�]\�����e\g����KIj�.~��*��_i�8�	�DH��Ӣ2Ԏ�<[���� �Y���k�45&0*� c�������ptۭ��p�Z7�R`�,)�[�H?U�m��uQUi؞p_���^���P�ħ�$����8�X$�q���I�_	��t�=V�z��8�>ٟ���v��i��ދ�3👩�:%0�]�V����{��DiԙR��t'X�_n3\�K�K��e�ܞk�3j���RX��U�TK=�������Cx��* �z�!$�l���|ZI�b[���\��$��[m�2Ex�0�;��E߇�t��O�I�f�v�דh��М���Y�� ��˗	��*�V5��hkީ X�=M;�/��/�9 �0 �`�B�`Tr�l��_|C�JucD��av���D�	���i0�eT�������z^­P�lNF�5h�s���|랔�4yhl�Jld9:�(G�H�=�ǧ�xmna/ [���i)甈���j��`����4��m��U�'�l�.�&��To���W[C��2��"��ӧ2�:26
��"�6s	=�ǕJ����5���z���K�|�B�N�$��=�CЧ��sܜ�Ǔ{�qo-������osJ���1�{�-��"�w��r�/�E`5\�<�$C��%�o�R�pf
+�I���@������մrl���N�*`'-Aӯ�.H;�l�%8A:/�
(�l�ZKV%��։N�!>� $���(����Y�
g�-������=g܌�)�̬�ʛ��F��ڎ�O����^fˑ�1���W�BΌm�{\㉝��8���l��.�������05��g�T���]zكH\DY�X�M��_U20Q
���t�mn�=p��xD�h����!;U�!�c���F�h�']��A���Wp ����P��A�kA�c�����s5~�W�kO\���A�\|�\��(T,�^��߮��T����%2+q�o�׉�����v��HENW����F�����:Dɩ���M��.����b����J�����L�X�),m+U���Z�\�7;���e�
�Y
�J�aDDu=��P�r�S��H&Y�-�8�V�]ʑ�`��l{�.���5
2�$�@��x`q��m��x$K\�C7�}BiV���{8jw(��<.�N��D�劥u�#,/� :\�]*�fP4?�����~?���Jb�f��8�'�d����~C���C��7�˴�x��|��a%������N�CE�c�pِ i3�~@P���/���}&�j&ZȻy�
�hF��ⱂW���:��*7�/���Ϭ<�W�2�M�,�҆��+,���۽Fysk:4�!G�����ܮ��Q��ٸ��n�*��n>	k�)�[ԚL�����9���;1��������PRa���WF��t,��E����B����B��@�����$\>x�f����a���K�q��)*�����7^D�!~���^TU���Zϣ�Mh9hW���J�%�E������*���O��8��S��r>H����r�$6��;��P�b+ְ��x�z�ն>���۾�]F�����H�h�v{ .�U�W�b��`��k[��]�p�