XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Ȝ&Af&�=H�u�`�J݌���TKk�J���,x�q���
��rR���hXwt�Ph(��]q�ތ��P��[��#
w����Z����ϫ�����d=Ht�	Y�|���T[��D�%<-�C∬��%u[H��V���a�lO��x������j����ǋ:�ȓ�yz֗��Lo�HW�a���yk>ϝ�F[!Ժxh� B������Y�{�c��E-�1�����Ī��p�W��}��4>0��J���!o+���}̣�,]2s�I��,�l$�+��{.�s1ܡh�&U�7�ü�̗FƜf����rԱ�a񠇄�
o{rz2P�(��{q�� �w�<��	�"}<�������Q� �G�$cHd������P���9����-��T&�9��)����f��b�d�Z !�C����t[�7E�5�l�/��61x�co_�"R����)BKY�8E�B��ܷ�o�-=(�cARͪ/��d���t6
��<Zq��}Q �:�07�ڽ��qM1������(�w]L^�Fmc��S͘����~Ч��(�9�C�ݝ_�
z$��&}�Ҫ0���wie����IC��`�X<r�f���/aH@�h\��JX�-��Ņ^g�*gz]��'L������3OKv�M���#uq��}�ea��|~יF\��Hþ�(7���ds�(2C��Z]��S��j�����*��MX�Vg��&L�e��e���J]�XlxVHYEB    fa00    28807�d�-�3����8�g�A���R­{Z�&,؏l5�I#P�Ii���z�M���%�w��Z5��	?S�Y���Ӄh^=���+�,6+}��Abf�D�R��1�+2cή�v���i�U�ѮaXd��ՆD�EJ�<q��� ��_��-���(�Ya�i�Z�;Wb�n�,M��d�
*)W�d2R��L�"�[J��ӈ���I��.�`#DO!��h3�cW36�A+$uB7�.,I�`�Ô��%}�&�ߔ�;�(�X^boC��yՖ
5`P����W�J���Vk��23c
��f�mL�g	4vZ$��ZIS��q��$X�Y��-ż�����|�[Xr���6d�j���	����C'�� �n��; �&�Gȗt�7����@2�j���>/1�D�m���ܱ��|��	�b��9!�D�)R6�Y�eܣ�tv�f �����T 	7�<���`L�D �֌�y�(�>Ķ�\�˛��(�j���*��1����'���1�1�&u�!�"���z��ۆ�[�����_{hf�pz`{��67����F�Is	�� �K搖`4��z�g��7&^)�F$f���4�2<:S���
�p�ԉ8i��
Ȍ�	���k�<� ��p������T>���Z����b��z��L��:�`V���E�29�2!ف!P�YV�V7�
���Y�zݜ��^d0�٧���;, x:�	��]P���zU���gY���s�sV&�Z�	4�&;~��-������G��Iwڏ�2�p���*�$BIh�(�;);�>s;z*���u�P-�ܑ�t[�d�g]��A(F�q�'3�) S��[)��olZ"?�j/	79V����H@�(9�޿v�u��ꃽ��� �¥X4չ�ju�3�fd�l¿���0��t�����"A�g֒��hpy|#,�V���9ϽA�G��=1#OsB�]}^�R�0�Q+	]�3���.̻�܉����+C��t߿O�յGM��,��B�LnR��:!F�u���z�G#~����Txwf�)z�1��s��2O�ĉ&�z����
S�y_�u��.K�����׌>��F�v�I-ʕ�F}V�	�;���'�����:����������:�+��%���m,�a	j�Ҹ���΋n�&�,@J�^�J�V(�[��^�����"ݑ��[������k�9�L�TJU�-ы�/"I�=�ߴ�0c��m�H��x�c��#v�~�>n�0�D���r%������k�oB�Z�`���1p*E4�s�s{3u$����[���:�g��[�:د��V��9��Tb�?:��5�$�{����.X������;D�F����.��.������9�pJTO!���?��,�	�~�;ŋ� r%�&���)����ێ%?f�1�׿�9xo���!^ݡӾw�F"�G�F� .޾��I�˨jei���k�%��a�����@�����u	#��%�a�{,�Fd�{a&�Y�ܺ%�!-��aӱ���#z�3�E��ݞ�� �3i����t�h�c9E*x���q�C�1�!�%W�����H�ch�HN8r�A�,.�i��%e|�T�(P�Jl��_(�a��;���D���������'e	��.�(Շ�pp��V�ӯ�M�Ky�U�׊a���"�oN$�S!�� ��/�hd��Ї��3��E4�i��X�� �1������8t��q6�&z�%F���bm��Phrŭ����bq�bZ��Q��F\`z���H���q�K����;���ފ@��3�n:�ZSՅXJ��u��/���KR���]�e�y�
��[M ���#�e����B4����O�_|�=���.�m�W*�sG�����@L��7�d6��to�߀�U�>쯍��Kc�����'���}=�ֹ�"{~�7��u��D��ț�ȃ�Bg�(g�$��C[���NI�&�9�O�(32���D�J!Sk�UU�=��D�����MS��\".�l�m�G<y�.�Y��(e�t,���iTyƫq\'�W�7%��Oڈ0���ЎM(�>����g�_V�,K3��U��NP ��D������]���0�臿�9`u�*TAqmV/���l���D�ō�ƵXS(�=Q���y�б����Š�<lx�h �#�i�ŏY3-�3<㨺4���3��Čo(�$)N=���Zr3�����䗚���8�Ċ�0��@l&Ø��D�
~҆2��]ɱس��e��D���4b^������^����"@lB*��������Rxч�dH��u@6F�m�����d�M.����<��ӁvӢ<����1៯j74�w:wW�\��a�h�����U�&Ks(�,�A_�sͽ���K��bb�]�ghS��!���P}�4�ǰ�Θ� _�(-L�SY"�ݙ肛�u�̆��{j!`���ڡfʂ�-�7���aOXS|��@�|�ނ�|ѵ�2]u�VF z�R����(O��A��P��ϭt@����!�fM�#"M:!�";-(q�7�� F��6��i,�c?�2p�oᇥ��r@�!�� $��#����{R'��Ps����⵪��d'i�� �F�2��YM�Z�ڝ�E@�	�9<8N�a֙V��Hx����vَ�Y�r"L{�>�~OTM�c{qG�M��-{ѥ-�ҫz9Dd�V�C�Y��	xZ���.�qQ�X�2��E�u�z�W���e$����gQ�/9�ǪN�2�pP���[�VF��C���>0���E}ʋ�C��^c����\&~X��U�J�8x��7�����xb~�M����-����yКO֝�)�+���F���Aw��\��ん}�@�x���@��2�%bx�>ǰCM���Gx`�	w)e�@��Nk8~݋\4���)�#��uv}&�6��R���ւ皢��,4g�
%r&S����Lp7t�yI�;z�K8ɖ�.V��(g�= OJ��q�ϒD[§�q���81�����l��%�◧�^v\�y�:�e���1�L�[���?>غ<V,|�Yf��G,/�oFz��F��K�O5Ï�w�0�/�ؑ�M��Ԩn�����&���[f���r����2���GDL���q�L��`v����O�,��H��������υ�!�u����j%T��wvO�Q�?���B�7L/�DM7�xfw��XJ]���ʅ�������8�s�]����t�^���n���Ӧ��>��!D|�4��5r���4�������Gd���T��{��8-	J���U�tE�	Dt��D[���Ш���(�i���ӳ��pt/^1���"kS��7��@���k{P)?�x�������9�K���g�tk�]��g~�j�51Ch��\t��R�vRڏ^��H��R�(��9�c2l#�`dg»�h2��� ��2ǫ�'�Ǟ�)�áR�gc��I�J�|�`�2�q�"���\-w�;�P�CZ��<g�a {ԕa��[�b����㿧<3�/W&�ɥ߃�����:)� ���Zʢ!���#�� u�]w�C|�#��;<SN�%c 3I�����]v���D�_��㮟�*%[j�� ��.�WP�)�Zx��:�c�ꤕ0t+�Y�D�]:�1@�'�N]���px�|���\��$�2������a\T^H�n�w�I�����3:�NQN�2�1���ar3�<�w�Ў�} �C߷~�\��X;Lkλ�"r �S2�4�	��%�Z"u��YC�������c�Q�l�F���@�gR2��y���u�5ȚY��~��7i�'Z�%�9�S6�w��������ڧ�F��j���)N��e���h1�.�9BNt�y1��.���I�C���[��v�ݜ��E|��opX��NGQ�w���mɯX"�^S��N��Ik'旷iE-��3����	CP��o�2�[A�,��g�%8W��:����{��;�q�Y���UP�|9�]o�?�_�� ׺����)9�̝ޓ!�Jt4|�%������B�j�A����B���7EU�P��	d��Y'��t��p4��W���N�)/��7d�8z5V�����|�Qÿ�-9R�����/LT��׾����[T�|��Sq17�\ٛ�P9��1Ku��x�A`�F�r�X��u<�w����"�ւ�a�}c�6�Y���X8�#�t位�䎦���-�bfEɹIet�I�.k�7d�g��!�~���eI�w�W�����X����b�c�3t9N���Q7���c�B6�m�U'�#6���Xb��N�W?J����l4'��G����ĥ�.-�ȟ�❝�����	4��]f ����Ol�Y�`���K�x��u 6���7ƌ?"��N�X���e ?ĸ�)�t+�X���%A,�� {��L�� I���T���d
o���ak ��9�^�|_��x��;��c_O<�Wl���{�&���^�����+��j^��9���}n(oHa�i���w��D�Zމ��qNSp,��G?�f��l�����2d���Fق�]W�~ǔ��zľ�0Ȩ=��� ���\g+L�=̓xH�o�Q�h��6�qG+���``;H\��^`>.��Ӈ\�����#y��]%�	��r��R�Q�l1z�o�V�L�K�����W���X�컋�ĭ���e�cGW�M���">�:t�bY�Y��Ͱ�HFpt��+vpi˴^T< �$\XW� ������׬��w6ⳮaJ�� 1<>���G�J9�F/��M���躚!���f������ҧ���#.�;D��HX �xg�<�I�;������*���2n�h.�������~,/C��#�U���ߔ�\o��������"l뤓7�:iO�s%��B���4�Ϙ��'3�M���_>���I���R��r����.���Fc�Fk��"c:��#�rp�k!r��Zp?�!P�*k��$!DT���������#TZ�8�1+�+�t���7	�� �Nj�X۟�J�� �\�]�.vhg�螅B@\JvX��Ui�W�2A	�I|�3�g�Ve���Zǒ�ceG圎��>�K�Ti�mB�����G\�Ϡ�h����G�% u�5��?H���G�<YF8��2�Q�.�����͉����,�G_%��y.,��4{z�xb��͞&���jɗxa[�ƫ�\�,�	���lȟ:H���رd�o�a���C��QJ[X/�s������F
�D��.bS�G/v��o"c'�T5�d�
Yb�1����X�5�����W_gB��]��\��cT��19�C�b;��I�X�(�ck�y��6t��)��k���������X�%8��3V��)�,đ̢g��Gs�:����z��䭬%w[����C\6"�}\��^͘˚{K���Q�K/�Z<��������@9��k�T����x����K�}㔪�!>��d}faP;�=�X8QCM���;s�HR��/�Uc)�j���\8�%������n��O����|,�o:����P��7�=F���LH�~�[��f+� �!��_��Pq��y���d |�����@�U��j,Qx��*���8��ŝw� �U�c�U&�v{c�d�0I8 ETkKj�K��$�|�1"2��V�v����EH!+}T	Bܶ�ht�4e`v�`g�5@��i"(8�HC9�i8��[X���Zq$�F�A��o��:���9��Nl8TP��Ȕ6�3��pw��	"<�$�s�]�DD&(�_�"�!]%B��g�7yO�u��8��|�r��J��E�!(�2gn[a,	7�g+����T�?:~/�~��7���i~"#C^g?����g������խ����	��9Q��Y�U*Vs��b"D��ECcVF��!��F�!���W6W��u�v�g�Y@	S(̙}cnVby��R�Y8�#�M�{"��@��'�F\}�.�Z_�`��RP�&�=�@<��;K�-���{�c�D�^�e��8C��}��OPô���6r�SP
�AY�籑MCz/�X	 .�"N q������M�A�?��鳖+| j�6(x��`4�$}���קͲUC��?���z��%�ہ�r�NM#�K�h�oo�q��,����t}�M��aa�M���G~��ً��
��;�ѓM�S{T �j�L��n��v{�'xruY�N6Uzi#h�<�44���-n?����9ޑh�C���ps 4a9�$fY�ҁG��9�6��>�NU�Fbm!n������ψ����lQ��8�SI՛�#X����w�u���	������ވ�b�Yq����',�!S[I=�ual45�e�D)쾖(Xl�=A����4���Pָl�3�H�F"?�)iw4C��L~��9�:mv[�W�:p����M�V/A�O\F�~�x���� ��8j﷙�->�E䟽�Wz�u�Q¡\�� ��-�c쥦qF��`���@b�P$d)�e/�(��&]��v���(U0�����`�=���[6^e����e�N���H ��#+\Q����~%-��9IN2i;������ٲ�@ړ�v7��d��>F���E�oe%�A��z�~�V���k[:�]�e������y�E�q���3TBw�w3u��T#7vS�9��-w�}s����	j��F� ������u�k)�IY¢�꿓�?(�0�n8����ϳ^7zS��1�
ހ�óD�o����M���1�c�F��������K���Ls��ɒI���s0��9�u���3P'�1U�MŲe��O��̽a�7�h6���;H�����*�=֮�01�}��v��|�I�����Y��r�9U�������'<�q<,(�Vw�<��@ ǦI�&�|.��]�/�K~���s1!�����WMp'>a$]E�_��A�E�O�G�E�Wyr��QH�����˸9�=��2�u�T�]D�N3đ�j�*��ʂ���M��'���-�x �<n8g��Y3��SX����_d6��ڊ��t\n�AE	�?[�M���[?��bg�*x:Z���?�Y�D�N��&��	�wJ5B�I��W�N�җ����Z]��soQjAw�7�ю��*�����BO ,S�� 50�Ȣ��[� j�4��K��}{�BF�f�{|]��?� ��0]�AȒhMm}�?���BʔCM3�:c��̛�m>%xЗ
��S�X��v�FzŬ���W�\}�D̕�8�[����UJzöR��+R��xx�0(����2� 
��9�,~�*A.��x����K�Y�t�)�ᵕ|nnt=5ᎅ y%y�L�^�s�o�� +ec����}���:K�9� b���O?��a�ѱ���ty��Qp����m���6fQAK?3��6b�qsl?���i��r��O���U���̦Qr�n��~8�Z�n;��!�P'��-.0���?�|FeR��_ 4
+E��Ύ�C�t�����n
�l�ex.�Ԏ��)Ǻ�idio<V�%��ѹe���7Ջ#e��\�_|_����L9��9P1��طy܈��m���)�Ik#Z�*�?�����*�% ڥcϊ>�;T3�<E��'�=��/�B�b"�DP��Sĝ4:�J�Ô���>��釄.x�P�O�&ig&R~�c�9���h��i���l�,R$s\S����!X�H囷c�F%����F_*E�(u�Sb*��w�;7�~�̀*�Ʌ(���{�~_�_�0آ�~9'���ԇ$���J:�;�RX�7�}�j�|�Zw� ��$��_���������������a�\��0q��wM��Q��N˪�����Q��:�,ïf��DdL^�}~��C�������8�W!��X6)A��t}rq�N~��yBw�ixA��bgWP�&�$c��P��ڙN��(�NOJ�w���#G�3�㛋��'!A`�`i>B��0 ,�	b5[�Y�l��s�D�������������_&�}<��F`Cx��2�iU�dM��C��K0Yš �}� n���ev]5d���7U��ƍ�ۃ!\'�	ɼ�EQ���g�6$��?7B^�O����*��%��#�\�(��w_�̩&^���5�z�uQU��5''�z<�h���{�0ʓ|�dO!��Ob���:�ר�	���*w����n�[��j�/E7�X�iJƉ�$������D����gxc��]?H��"S�׮hU9m�b��۲�(j	N��#nS��n����
�}7\�!� DG]@I��+%��G�����e6��ï��PO�Ȉ��0շ؛sѕ�]C����r ��c�v6���,�跢͉���r�]������]����S!�
d�)��ƭ� T'��p�c�Lf�3zC��2���T�5��k�ɢ\`q�A�z�.1N�$ٮ��	�Zt�8�'w���H�h�����9C�7��Ez��pΪ_�?- �	d�Z��ߕ����.zw�Q��[<k���4He�&h� z-أ���<��޶���
,N���(�(U\�o8?��9~	���۰>@��xw�����LQ�>�w'�g�z�tC��[�|�]8����D�Ip'_�N/��P�R'qP��ˡ�CGu���-Cs@g�gG�7ԑ�[_Sd�	l�aQ\��bTW��e{K�����ڌb5f`��͈���b����]���J�Lĥn�A8��Y��ت�{ڡ��k-�~��"�4p�ފQn��B�v>泉 q�|BVѾUU*��v�7�&���?$>d�>���A���]D^�X�>���禑���x("��\U1��o�M���i���H��r'�9t���4
�i�<7����� Q�ҴoQ�^�0dD^;���I\!s0`3�t:)[��tgł `||���0,ڔ�7R�:d��Ծ�,��nj{W>ZG{��Lo�!�a�.��[�h
�X���{,v��ed�d��
#���Z\-U����䬗�L��t,�Tr�mr���5����4ؘ�^�d�T���~�;h��t5-��2�7�f��߆�mԘ����ף��\��	`T=�D��'�T7�%�7��3���Z�G�>���܏�j&���ѱU�h�D�0x�����:1X���>��*��{��h`f 
oifr/�a�ԇ��ս�r.`�S�w��3��p��5��NP5RS�R�?P:�(Y�x|�b��Ï�����!�����4�ne=��\��ꘙ#�%iӢ�t�#� �}�t��V}A���ű�7-����?G���;▁�-�i6f�� >4j���l�՟c0Z4�~oJD!� .�<���v�5���Ze3����C����hZ�J�k���J�f<	P�ƅˑԪ��4�|f��{�,1�?�}O>
����iד8 U���\� ��ڏ;�,��� a������9n����ak*�\���=�^��n�?�#��qk��i��Lw��U��]#��5�<Cn
�����Y�e�� ئ���������>|���c[�\�J������b�G�C�Q��D�6��������v*��w������U������2�k �͙u��?G`�sH�#^�]��Y��'�,���x�o=���CK.��^���ۭ
<��q	4��)���/#����$:�KѾ[��I%��HSDA+�CQ��T��3u�Q�n�MD�X�S��>�!��ZJ{y'*�"���]�c���F�yL.�m���;tN�8DQ��@�+�\��:hԳ&~�n�=�!S4�1y뚥M�!�C��	�����=Yg`��8⮛��0Զlʕ�N��,�d�?��A�4�RíS�#��7��1� �J���hd�T%Q:?_.q,1��jM�VM�<g�!�~�0}�0\�l��u��~2�%VTSOb��&M��t��V�1�l�>���f4Ξ��%{r~���	/�����X�����P�`����Iʲ��gr�έ����-�x�r|t��&�q��X��N�7��eQnf����a�� �V��Pp�d���Q9�D��b����9�Ƶ�\:�}Ƃ�3�A9q;��:	��v��x���?OԈ�����M4sLG�gCb��3z�)v���ͤ���z�NEY7{���X`��%A0B������7N���XlxVHYEB    761f    15b0L�W�M%��[7����B�����zOޔZ�S/�%ׅ�T�G������;�_H{R�I�UB<k�D	�5!�����#�
�\]dK���L,5�Pn���	�g�;rl'��Gϳ�Mta\�����`��q܃��]��G,S�����~���(ҍ9sَn�bP=kP��
�ګa�����ю� ��#��M<���N#3�ew������*Y��]۹�	��ۻY��W�����ΜO�S;G�Q��g,1�a�ABg�p	�sx�4^h�)��b(�X���dFT�t�3��l��8M�V�����������L����e~��ޜ|�P�)=rÐ?Xp�fs��͞녾�.�;�}K�u��[+�B���03�UC,��d�x�z��\V0�]��lڅX'5������ �ݪ�����o������tkw�V���J����L�Hƈ��$�%�L�.�''�~�����)�thfC��!+����\U����`%~������8�\���̲�>F�brqj���Y��
�r�h|�:�O�I3� F�K��ñ������-����͠^�����c���;�D\lb۳��t�	�G���`�s�O}O|e�T��0`cs�\�'{f���v��΅�A	��񸟢��Sꮿ:�Bӟ�ݶ=�a-�d�~�.�_����/}g��v�$c�>	���m��~f�hΗ7{��[�uK��W��@�`*�^J�;ͷ��A0'�`a0̇��:۰ch����[�
��Me =�]oS���Ӽ������x�1 ��_� 3����B��I�᭵�R=�)s<J\��E�"����ξ.Q�mk����/�d�o��!�~t�щ��A���X����0�V�W�M�*7@��>���A��������)j��m�(Q&鹈�*o��4.�n�g�Z�$�w��)�w�x��0���M.`R���F����R:�9ڸI6���yFa9��u��w�+��\}	?�ߐI�t$�B�L�H�T�1|�#Uo �i6Jp%�����8r6zg�s��9��U��|@;�~g���qչ'K��љ���©���W�����4��{�|��؝Ǣv%.Z�5�D�u����hw]�9EF������I<�B+�p��X��r��QT&���Йg�c�jT+(7Z�P6YuA����B�W�{�~�5�%I܃5kx������**���^N"�"r���r&���o�lQ`l	����SOO�Ad��*��PzW���<AV��h�¹���|�&��L"�M��n����DH�@����ۋ�~ı�)��p�=pׯ=�Ka;g`�b�?Xx�sY-��ĳL�$�4�ٳh\'��g���čA�m����u�?��/��gv{h=�""bUk9L�I�����~"{,s��t�Iy	!7�����0<�n�j���_$;�JDzf��*����p�v=����OR�x6&N�K-:�����g�N�$1�5���5ʳ<r���pk'���(����5%�}�G퍤�W�������-���>0�y׬������m�'�౻�2�K�������y�BW���x:eoYkù+�~�kDj�w��<}�E��r��za�j��9�j�4�@H����X��%��"%�I�L�y�ʑH�������7��e�_���P�7\A�Ʀ�м�4���N4��琮���
�,�$���N��D�ߠ�~ R�jn�O~�R׺�Q��qחq*LE�>Dz�EZ,��c�r���^�I��� v������1�"�y����N=�:)�R��5��!�D\����.(>�MP/�v�^���O���%�d�O{��OʒA�~��Ǳ��[R4��d99�`�>�$�{�$�`�W/	�ѵI8@�	�J�f/9���+R��~��(�zU��pi�M�����R!�Ƀ��d1Ȃ���ӿ�Q�uV��|^����DM֙�w�];
~>a*����iT�� ~&B{�W��%��ou!�:��}��p	��Q�_��4J�|'�w�������`J�������9j|aivP��;&{�E��{W�,֎�RJ������<e��,D���e���4Y-\剷�4�c�>5�%mC�^� ��l��ؑ?���~����>q�&������nd�o�)��*u}V��1�e0$]L��J����nȹ��0]k���  ���{񩘚QX�,Z��3'�b�-����.�Oo?l���?�X8E���1��S���W�=��1�ZG�ޯ�ӕ���[��c�3Mto7�����:G~~�p� ������ۏ�]��Q˳���y 0�t��:���\ۀ�������o��=���]ϸ"I���kU�h���lB�y�#�<D���Q�n*�=x}������`Ld�%����>r��Ȇt�
7P���K�-� E?��DS�T����9%ɬ������F��|��,�[Z2��b v3����
NX�YyDBZ�f��E���Rd�l�C�&��)�&|�����v=��!�K	-�����"@���y��H�ٱN�&K�����@�p�c��0ɢ�G��0�_�����������Ŷ�%�*��ޥ��r]O��Ia�\8�LH��Y��x��cY�[>�����JlR�I���ԍM-s�{����ej�VnW�rwFG�u�M�����(�>��ƭ>�d�PkA�uh�ެ@�[�D@$�6wr�Y }F���� +��ÎI4�2�����}���!�ޞ^�(���O�x�� ���K<}�Be� k~��P>*сP%���=�$�'h�gQ���=�C	<��·i�K��Xfo^;�4w��e��ΑƼ�R�S��fD�\z��a��+���(�ej�R��������&>�\��?|4�����z7���5(����[�1�gm�����l����(���yy��#\~�Q�L&l\,�酦d�U:���1LkEr��h��w��x*ɧa_�;�����'	��(�udN(Rg��v�/Ϩ��¢��.5��Ev��<���➂K@P��W�h����{o��|o{I�Vc�5=��\9sS�O����6��H�b�@��v��xԵ�#y����@� �FS�0UT���Sy�M��!Cs�?fzf/�a_�0�R�[��޼,�B�@�,j�с�q�һ� Vi�t�E�^��)eݯ9fv���џ�n��1���}e����:��$A3Ȯ�p��C�T�������eA�W2����A2�e��S��5ԝ�
)�T%�
JU���k=>��ꏴ��$� �Tƒ���o���Ms�}:^WL����>���[��HҔ��C'J�h��VƋ8�0y�F�V������-zӳ�pO:�0?���s	�U�?2y�]ASi��9����Ф�Ɉۤ�8����G�k]���Q=��D��˔}7χ�m&��R�f�T�U�*��W��Sv�ż��z9U'��Nt�	�,�ć��Y7z��NjE#q�n�	���z�W�l���������ѡ�+ՠ�t(Q��_ �,j3�[Kw�9K�����؟J*���[,�'�5hKB��۱���7���܇c���p� =���'�G#��%ь�Ȕ*c���S6�yh/G�mi�.p�F~������a�J*#}��Dip����.QwJ��� �G;t�P1w&�'$ё'Hva���~4L����#�]�lZ(�	Y�jb�Lud����k����M %��e9�V�hϺ�B�ĚaR��I�	M���$)_�\LE���~����9�C(+U�jiy�G �Q
��x�6d6�c3�c�&]3����� �H�;[��j���[�fkYD+ �`+��6y���e#���;�w�x�����ٮ��n��=���� ^��q�~�o��l<�����$��n��qb�L�{���W�I�qt���'���ƥDnX�j�e�*V&nM �9M�e�u����(QA��:J�!g���/m}��П9�k����͇��,��s�\q0l��(�?~�{�%�8�c��:�%�ʱ�xs�0lI)�,]��K�2�zp��ݤ��F�UM�O`Evh-q�uD��t�w��8<f6K�K,�gr.��,�{0��I+=k<x,І��ڹ�I�:M���2@Q?�T��1|(*��pUO�.V��SPeb �I��-�+�q
�e".�O��?m�|���w���b��1k����8Q~�$��g� �V�1��Z�\z�����AvZB���7��P!�=�a��<��JI��;i=0n"�`�=C��ܫH�{�C�0�U	E'�/qt�ϒ\��CzJr������&�k��6LEu��d_�z�'�6�"��3f�â�5����b�����[I�+�R��G�`�2�+��^�?��r���
�B��t��JM7D�eꀺdDi�|��0�щ"-���*���Y��#���p9�*K(Fj	��\����[�l�E��;�ޯ����20���D��*tyϮޫ(ß��m<���e{LV
䇦N|�`��o���Ƞ��7)B"�s��][������@[�гF�����=��|.�\��ӊ��΀ t�8��1�V"�^��!��e{�ƥ�t��.�X�^<�&��� �^&���汷'qc�r�Ӏ�	N(��ASz�jl�:XZaP+��s��a��W�4N�)�c���!&<'Vn}����<���Ƒ<�o����I�	Z�"���=��-4��.�R}�����u�4���߶(Z�� ������� ��W�Gwz[���̓����v(��  �Uꅈ�2|��h�l&��	"0�r��r�K�+l	�� ���Zp�$r�;=;4dB�[s��+h��*֣�e������5�-�Oچ�W2�#�c[>%��Eӯ�M��(��0!�ICъ���,7�󬰌x"����I�_�; [�YD��s�m�RJ)̒�L��w��&0���� �DJpC(�������2�{��#�<���¨��U^����$��ˢ��h{a=`���s}Vҽ���X�t���t0��46(u&��Rk�b�����.�Z�Peų�$��-7��� �͝D1t�:�B!�Ѱ����%S|��b6�kn���,�{��Q�vz5�:�s��&Q5��+1�ra�N"��"_���R�)�%�C£�ڽ���6���g+o�sV
V�鬍������P��i\���~���"N�A�w����D�W'����g��-����D�
�%���^k�1)IW���;�>�$>�"��g�'d8s���ud���WÛ7����ǹ�
V����2�|�"���.�r�J�^��[1��xx�e���*>�rz$ts��������^Q����F�N�&���nv��,4���5��t��sB����[�Kȣk7�[ny��*���Mݵ�~�C����t��