XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���"�F�dz*��
%6/� H��Hs.��r�P������5L��kN+�� �j�Z�Z���0�������� ����	b���v��z��kO��N1Zs%+D��P��j0&%�m� � l�7�+~�a!{�zj��R�����|j��2ݾ����p¿f�/��"��� ��f�mJ���/:�ᴷ���m��%O�蜜���
L�+�[BǤ>lfWԿV�� ��������o�t!۰�a�KR`�u�T��m6�Ta�bz�"�W�;옵�@q��p���$�������>�>Uc��������0?ɾ���;
"v�7�]��L?��nF��|��p�U]y����h�����J�:S��~~gy��J�r0�׍G�	--�i�Qj 2t^}��[B�kah���S����6��8�%M�9G��r��&�'�݌s'}�ӿ�1C�t��t��B��k��ze���y=����a ���#o!*l�����>�)}�YJT�
�R���7�C��ߛ���eEɚ,(�u�	��-d��SIBT�{׷� 4��ˣa|�՝ٓ\D꣥KQܳF�W?�ꚳ: +u���y����=��"̐� �l�wt�!�AY_�M��6� ��GX/۽m��	��Lg&(�R�=���z��?s�W��4��[�Ƣ�R��`��(>�9��1�8�@o��аA�d�n��J�v���u���?�E���/�,����������8�<�XlxVHYEB    4a7d    1090�����'eX�\M���%���堢r�v��*W=��� ��Ě�sB�"�(��4MXtM��tv��țW9׃z��t�~_��������h��������w4#YǏ����>�*aR��8�Q�P����O�v~˵�����'�_���>��1�gdt=~�F����hnv/4�"�su^��1�CyGĹ�q6#Z�J���*���d�j���+���n�j9\�X��G�$,(��Pp�l'@id �����B����./�U��͋}��J::��Nd�����:�C��� ���Ýx�2��E�1Q��6���NR,�R�}�R�����f��-�~�C$g8�TrwB<��꽟���gC��>�葝�2b!7�~��v���Q���u��"�Hh6+2n~�@!ko���o�<"�(F֎��rr���'�cs|��Ԟ�s �NN��?%�]Vx�I�*�sU�~��p���y��������Г�y��5p�yf¥xd-�=;��Q��8�� 'KT��1�𑗉�F�p��d���8��2�w��,�E�G�q}��Cd�}�9���Wc-�q��l��e�l�����G[�\��ϙ���p떛hf:̪���� �&����	������h�D�xh؂��!'3`8qQZ�ȴm��LN�Xn��l��A����K�Ϣ�7*�l/�ܖHH:ȧ�$��䦂Uģ�L��Ќ߆of a�7�莝=_[,��J�h+�?R��vĶ����VA:ЈT����B}�x^��=�?�1,b��a��nv���)�PV�h̦��`	Tw� �ߌ��A�5��[���+�U�Q��|j�|	XF����%���ZL�A�T^��<�O��q��gn8�f$�Ax���в��V���J�m#�X���WT�Ҏ0�ƪҕ�ηvï߶��+��%yz�僭tG��5H����8 G
$CV,����X�ז3��#���4-U�?��6I~o��М=n�ߛ��	jc�w��a]�L��-�^��ik�s������i���u�������4�!<��)�Ge���!����Fc�{�A��=�SE~�{MZ0w������0be-*:�Bb�Y�A��W"?S��͈H����qCaG�,t��x_���c�7�����l.���"*�rvR�M'��^dR�[�} :.�g�o������0���1�fz;� q�6\vbKy�!�$ �ɪZ ���_��RZ��۪�G��J����*P�G�yxw����۔I4��,UrR�(,c7�<l�I��_��+X]$�(o�m6�q�j�]�g����1@��"(��5���K�ڭ����Y��⏶�+�|E�,�t;�r��n�A/v�*(���_�!T����i JT�3f����b�2Rׇc�0�ل�9���Z2m�)[C�����)J0�}�B�TO C�����l��VTɦ�̈́5���Q�x��w�'��uyta盠�6�9l�s��܂m���������7[/Y�aEy�2v�Q��`(��h�����獔�ӟ��8՟��\��3W�K�	��	�~o�n�P~��!���ZՊ>Ǩ�����.�~3�����ܐ�s��W�w�.S)5=�
�4ynG��|���HI?(A!Pݯ��������q>8���1�ql\��Xƥ�m�UEv���fO�pa�-5�b�4� ;ꋁ��Pٓ��J^�cZ�� ����rd
C���T k+�P �sMݢc��$:!����<���z���m1��T�1f3��| q��R�FT���T@�]���Qh���nσ��C-8��Ik��t�򄥡�5l�[�D	�9�qW[��h��! p�	%�y#�-��*_d�*�����󢶞d�@j'h�r���h�����Em?�+:�PB�9��h���"g^�<��a7�~s O�%���&Ylc�xX=ji��űv��M?w���K��3T�[YP~n̰m8?�bʒ��M��Irο�J[�r�<d�5U�,[%�}�˥����1Z�	l�I�W�s��m#Z��ju��ߎ�DҾV�G��0�Mc��Pƶ���M��| k�jb��m=�h�i-��łVu1QB}����eِ
թ�c�n4#&����S�H1�t2^��ک�:�D�ci�ßq~�}�/1����:!c��؂���$������̦7�/�^F�ۖ�W�#x�%dM��Q
wK��E�c���_�9��j ϗ��fH�b�D�"bzS�T\pJ��0�K8O��`|�ٚ��jW�BE���p:H�צ3j鼚�:%�b�����M������U�V�����5qu^F�O�CQ`54B:��P�v޽D��T��b��!g:P}���	�Y#��V&��^y����5D��$�X�\�q����|�A���4d �w ?H�6b�{�6W1�1c�V�㲩�cHZ�_'�� ���W%��\��g����!A�쭂�r�lQeam��]���Ky�,�9C����I�Z�J�Y���Z=V�1����7��6%S.g2�|GL����`	�/�ŷ)Y�Z?\����;��r��O��r��՛�b��`���\s�D�.��Oթy� �{L@v�B)�O���f(���h�]3���y䇿�޳���O˵�)s����P������I���l^����pgaW�u��*˘AoC	��M��������^1����j����B��v�(���ƇO<��!3�M�EW��-4)�X�y��B5P�g#k��;�ex���r�-}��-ɕi9�X�p�&�(l�D;���m�Gnu�ሕ���ܯF�ٵ����R�-j�/.�!�oN��g�0�7�*��ˀ��,�FJq��T:�&D����a����䈽�°@�Ew�Vㄼe	�E��!����o�Ȋ�����)�\����Δ��Ζ����N�c�)u�)��Ӹ<V� .d4�	a�I)��ԯ�M"xt�4�m�DV��_��x� 휕5;( �#�����FU��,��%��q��7%�a%�+P���)$�?x�uOډ�-H���*.μZ���}W��N�X�k�L(�R<y� �G#�;-ƃp��c�\�)��[ʸ��9��,w�Wc� ���I*�Hcz�T��)ȣ����2�L�����{�A�z�����b�:���r��J�;��z��#l��+��mE�����1<SVK��n��fv�r�8�*��(��);ts�)��a�Wb��
{7�Ȃ(sη��M]��,���:�#����î`nŭ�����l[|����f��+���)�8 =8����V#m���)F�oO��pċ��K蝤��+(~K���ٓ@��d+U�~���
�bt	
�����/s<�E��@�Unsg��������Y���;S#�c�?e���G.��1�D^P�9�UA��ay�)M���z�ݎ�k�����w�(�s=i��| �`s��ER�����w���{n���*"�w�7�*i�7	lO��t��<W�>��涅&[z�I�C��C	�;�D�P|��\�Kv�j�*j^���{����������C����~
��M�^�EU�X�ot�dh�&��=�Z�w*�
u��KK2�yb��Ü0��F�X1{m絁�;������=�'���rJM��I�����#�$����$�SSF�\D�h��P?ӼNst:�J���d�w�?^�+����ɉGİ\6�?q4ϻEd�~�o�����S���� gn"�RB��CRM��rnqH������Ȕ-�cſ��k+����{h0��L��m�n���@�`�^��T����'2�)ˌ����χZ��<��/NI-��9=_���!rS�|���O�x��\�� ��x�`�b�;ί��Ց9˟��-�3;c�E#�	n@��ſe�X;N�h�/{	�H��X��1�^p����.3�Dw-�m+ˏ6�rrr56̏�^��heu�����|��esMR�S�xc3<�eo����"?��r�ڶ�F�pQv�e!�����Ƃ��B�2�خB���U���̄g���7�v���Z��ㅩ�{cP�${�ȯq�dM.�N�U"�۰4c��0�>�~��R�Cᜄ�����𹊿ObD%p����~]9bK�DYc�e�j�O(�%&