XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��D�E=���	��#i5t��
h��3���`&�)z�{i]�S��.�o����tm��z������r�^���D�'�R��:�$��=�g�=iWzƯ
��`j����z����%����W�J����ۡ�_�3��RdN�H��+�����"I��#Hf���҅�|~�Pc.���ep�[�Y ��<�5�^��K׶�!D����TO*�4r���)��ؤ�b��h@r!H��	�����+*��?�>�c���vה�ڹ���� ��?XF�p�V��
2������LB��uYp9�&��ԟ�t��E�$Il�#$cJArd��ǸOs����6�"�:�B�	5�[s�j_����9��	�����M!���k{BNg�;��H�v���m}N,v�q����/�KJ��H!�F�Eg����E��/5��;|�B�[��:N�<�j����4��~ޜ|�7�Jɬ���OQ<	��V�`L{kU����.����V9��M�3`[{���[Heg4K$ݮ*#�Q�b����2kX�vt�1��a���夡="�A/��@S݁'Kf��>�]�Z62��]bG~�=��:��.gM����_|͏ԧқ�n]�B��0��S_3�Uݒa�JwR�[dJ�� �o�2�+;��z<oPh�=�9���3,�/��]��h	G���ܶ�p!��Q��l�_W�|��2��,"Iz7���j��/��� z��+25�>�*�D�Υ�����]�����5��%a�'XlxVHYEB    fa00    2470���+E��t7�r'񆤸���sݗ��r�%"|YV�K�����8-��f����O�a��i? ��`l����G�x1-��J��I�yM�=�`>���9��y��|Mg/�)����ue>pW�DX~J�R��2\����@P>ҩ��G���6]�=��Q� ��HfWxrt�}ɔ��e"���X�>z�U�ݖ��m�k������Q�H૯d�c�o��@�@���2�*n���X�9��T�� ���f��=�͆�U���j������\9�O�y��C?8��zǀk�c�ᗮ��kL>��d�d�����)��L��md���e��@�w��F&Ƿ��䙔"����u�{���&,.���^�M�;��ҭ:�\ތ��"��J(̗ N��Z���=���+:��� �a��Y��a��?;㔫ݴ�[��k%&/��O�sL	��\ַ8���+׳�Eϋ�A��oH|��<�#�Q���>@`���&M]EbK�KH�ۣ�;�z��4*)Vt���x2IYJه&���c�Mc,8��=Ic���;��jQ9��%,�RR5�:j��d�)�[�lЁ�������i��;�y��'sv5C��cQ�´}Z��~g�{E�L��5�e�ypc^�����v[�ʹ�^�Y�1�~��Fx�C������L��' oy-^�g��+9�d{���Ao���hu��AA�{o*Җ� �%ET���8o|k�{���i���"�}�	{�}�������7#?rX�WzxV?rV��h��@�~�����9����un����^Y����u/c홉�������{]�,/#�»��_̨s�t�O��e5%��hj(�f�	��L��;}���������=Qw��7g`wnL�����.u�-���Q�,��gR��_�%Y����?�p/$T�73�pb�]Ta�R�󠄉�4S>f[`t��M���6Q<���~aة�a�]�Uw��y$u$�V��\�-��
&�l�ה6���*^�@:�W\Դ�2%�AF�X���eu�Ԑ��QU z��|*{����(�����.�L.6Qݜ�'x9��������$a��(�?�	=�1�2}��
�>�/2�$h^��W�'�+&_��	t�z��n��2nY�b�)���p�%TiD��@�1͎l���1���5*�����[E�T�Y�S�}%����=�Γ�Bv� ��}4�^�l�⎐�� WG�#~}��*��a/5i�z1ϐ�%�}@���]B�Z�lW�;���R��F3k�L������4,���-�Z�D��A���]BY]�o���CS�df u�UXtC�yk����#۸��;���P[a���3��%ܥ����O�6����IZ��\��8����n�KB���S�a}�;M��_/��\9ķ����B\�	\A���?e�ɲaEOE*B*mŹ��p�!v|ZJ���|[z��P$xQ_��C����:<����ԒM����]�����0��/?�b���� i��s��'K͚����a���s�]X ������s)|�$	��?3(y\�)�j����Z� ���G��Q�F�ߝk���}�\D:�
<������'�oQ�f�z��ڮF�i|U��� ��d�������v>���z���En�傚@&�J���k��O/3�[��26U
�}+L�y���>���K53����6Z�q��m��|QB.����_����}�t=o	X�>>
i�L}�W�\;�A꿽���n��Ѩ%�X�x*LC�6���L��!ޣп8V7-�=m#,3�ߣ� ����wFi�K�sYL�kw�02[LM?\v����i��"�iJ^���5H��y�YO�+���
-�j߂�~p)� b��*��91����t	ďn<!��h]@M���g����w����:��DWT��N����ڿ��,Z�4g�Ɛ~ȹU�$�m�,iO�G�z��`��
Y*VÞ�:κ��'��]ʸ1�~���W��P�5�,�X��[ElI�l� ���P�LveCY��QW3sU�b>�pL���:���@ߦ}�ez�|�1�K6�@�Z����7�S�V�i�@�n��$�g�e5���l�ɰ�`a����t)W� ��.:RO�� C�fmH��w�wLv�a(,Tdw�K"C ���A헬�VjƼ���Sx�Gt��M�b�`��'W[9�	��t��`�kR����>Q���%�ZQ�@T��Rd�S�J��ks:�P�.��kdu��о8�֫ח��3N�_*H[5��D�(���8�x�-?<��y���K���nd;�g��1������.l�L�1�aH���[�>� |O�'���¶�Y6Ä�j����bk�-5T>$F��3eg�*�7�H�`��a��9�f�j;]�!��2Q^'��/�Ơ_\i1+��M<��"�Xɗ����/��CnG1�Y��B?�tRS��r��P.�e-�%5��s�z�<���Ƨ��<o4��e��^��mUz��'�?��p�z�5iV�\
z� W�QJ/	�i"��⁢� [�F�٣�jf�bkQ�Rd7�W|\0hW�"�m�t7fq4&��?��#N��Yp�g�U�A��2w '��W3�ç����#4�k��n2�i?j�PH,bI�?uж�_a	��g$���r9��O�ʦn�é1�_�u�2��[6��KV0Q���D��`H)���t��w���7aʉ?TLZ�lw�G7cj���~K�&S�YR�9>:�a4�[ܤ_ �ˎTw��(3��p콢���I��쁂dh!�9j�C�`q.x��b#��x�Qy�Q�b[�"��
7��/����V�A�:�x�=��y��<��f�����K�������DӃ���fn���* ����.�d�pM���\��S4� ���9��̪v�����5̚�H���	879������%c�"��Ҝ����B�V�3
!ʩNX!�O��_��G#��"R��r��9������Nީ9n P9��}+�~@>U�#�D���
އ��F��>����C�S�����j0��3��I&��eR�"6N�Q�O��-���d��S���-��� ��؛� ?�ɯ��*�����P��S~Z�������L�����vRP/�N��r)@&H8
�����Z�h6� �ƾS����8�F�>ܽ�J�E����s �P�u۶��f��c~�QGYq�e~���ܑ&���ZO����x8��>��ܴ��:ĔǏBI����j�A�$)>
�G��C��ò�8?Lv>V�G������`%Uk.I�P6ep�ym���^.��83k����Ӣ��,�h��dr�����i���G�L`��-�D-��,W�lx$I����'1!a�L�%ȁ���N��M1[G�!�����F��/�끉/�q�ǜQbE��K�'���@��C�,����r��f������r\�Ѱ$�ʵ'T�@�s�ϟ&B�{�%�Ya�D��K�z�_�%��mA��v�+����r��$�◌O:̌����T	6�M%f�#=S�����C��^z��ő:/e�[���VQ*����C�in�c�_�$�g�����@\�,l�H��l��o��z�+��p:�vvByu͂����'Lȓ�K���uX0�l+oנ�K&� �������7[�η�+?񦸪�7���IS[�٤@�֣�̏rq+��Z�IH��)�'#�Ҟ7"wt��8I��w�Ģ���T0��"3�c`F4��_r.� #��WW$%xd�SL�;���Xg�{�E��5��A!M��ٞ�X�(�d����bƅyLKJ���S?,�B�
ƅ�r2p�\�ٟռB���K8&���8�D8�X�)n`µ>���S��M1Y��K`��DrqE�K+���/��]�(�Ղ�����K�$�z����maϡ�o�Ap��:h���gf�3��.�r��t%����@���Ɯ�؟Q�E�-���r��PǎE��k�h�i�{ey)3 �9��t83�9C�=ei7-=Jȝ���w$缢e2]�$C!�%x�S҇�\�h=hm����*�����W=��o�Zt�y5��ڤkm!��{ޱ*��3O����P0P� %t ��nwH}�.U	�)Z���@�1�f.��#���`l�.)^A�G\e6�,�ߩ4~��^����<aR
�ہ�� V��/pF��4�W�t��M6����wN�L�������%�9bu������_`#D�����
�2���tOb�-��pO���q�;��?���F��8P�N�mE��3��=��3U�	�/"� �=` ���)4�']h�9�?�8�%ߔ�jG�K&���4�'C� BB����n*��C}�#C3�&I?X��Ҽv],G�Yy�9}��;�����`�-A6 -N�P�T�1KJH�a ��sux\��Ǔ�����+4��m�[�r��-����6ɧK����/��m��E!����^Xt\1�svHb��#_����h)�C	�;u�u_�N>f6��k!G"iЫ��N$�fH��a&����,��/�ӭ��b��f��/wr��[�����>��[�H|1(E���cW�JR�y�W�� [��L�$�`j4�����:}�l!��x�����-���N��AJ�Q$-���e
X�W�=������{�G��.�3�����u��F�L��^�gGM�3j� E��"w����zo�U8����!���c,�*��~��,I �R"�_,��(��*�tb9-�r����H�^m��:H�z�����"���`�N3N�Ls��,�,�m��x$�+�����	�8�0<�	FH�nڢt�v�5��א	jSA����Q�V뙇Ղz�)�������z���}�f�[���߮�a�8(ज़X�h���֬	�����ռOop�r� A�f%�\rh�Fu����N��y� &������^Eo��^�xة��wKޝ�[�qR�3<�+�Pg�1���"����M$�E_QcE!�"[V�8I�2�����Ĳ䂐w:/K{~�M��(P���!�����+`ap¾��n�_�^�q�')�����E���a:��Þ�(L��f���*�,<�3Q��0:��!�Q-��#��4&�6�x/~q�5�P�A�ʂ=�4��cCo��������� �Q����K=?oY��^8LS@�/�dC��N�p�8�~���9qq����'��_��u�M��I��6���M-�Aq��e?P>!3�3�f��>�@�����7��&���y���Z���22.6V�"q*�{EF|���i�:5Φ�w���l1��5ӿ��f��H��ڜE�S����y�&s�p)���a�}�Ze#���6�Ĉa��Y��ˍU�g���[r3:���}%$+�=�Z��޲�L��`��%ǢXUu����@�L��^.%�'�{�^<(��F[x��������r�I,!�l����F6�H r��E<9���-�͜LZՖ�����<�ȥ�i7��S���a�/�p�bT�WE���3�|���]]�&d��^�z6��QfؕYd����0���Y Х]��Q9��IM������Y��� �݀�?+�1W�P2���kzq;���]��+Xa�ՙ�ux�S��/i�����W�榉�8�`�p{���y�Ǝ3`h��T������O�����<�E��nX��8�Qm�л�������Ni�ёK�A���8��1��j�Qn8&�^r"�c�<���ECqdeLN��� ����ܙ(yˑM�5ߒzQ�Iiŭ?��Z��<5^]��ON��(���|ގS^���c��ӗ�&@��ƛ%��\��99q.���>b�������T�t��#r:�Nr��o��rE�ᨨ����I*ʶ,�Υ	֤m(��D�Z�R�w���sk��I�m��1�0���8������,q��Ѵ����Ѹ��@G.;�=����"	��U�R
,��b�F�ޣO*��YC�K{�	ɐ�Fd��}Zh�ݾ�n���}N�GLʛ�`_�;*@44dNDc"�D�#H�{�q�Z�)T���Q�?5�C
'�P��6�Cf9�;�_%C=)�Y��dU����'��d���!N���E���bZ�qج�
i��z��ja0��u��m�ɘ]�᪡JT��)3p��R�;5,��ϙ�mE��s}1�>G����2+)�jV(�ڶY������I�B��������iƮ��ڪi�C�pj�
�P�@�d�y����A�f�4p!����Y�{ �|i��!� J� ��
�/8��V�� �z��L}�4�X��Ś<h�t���O��n��w���*��Zm�]��^��k��Xc�y���j&�d�j%*@�\�G�ӓ����B?�?R\ C���*�p@S2M�3DeS�� �b�g�Vg��	��`7'��g��*%I�T�>���!�@?uI�1g��4�]�5�>�u���1��Fi��i�� �>�br���{Xvj4�t��i6��5���N�p�)�͟G���{(69�xW�����>�Wh���ۿ�"����M$�K{�݅�H Րa�g'7��;�{�����Y ���3,jm2B��`��"�9+&�ѭ}��E|����dޖ��5�U������9�� 7g~v���w��lpFgז�k�ZQ�D!��=/��r/���/��q���}�4���Z- ڤi� �%E�},k���k���n��O�ݹ	aOU��y�T���z��m�a�vH�w|�W���>�PO��Yw1I�~5�ڙ$O锘&�)͏%��\����'v>��r8�G�΄�eEmy�8Y��&��ekZi٘Tf��5��H�^\����zNn,�ҍk��XR��o=� ��1@�=[pj"����96|;ƁH��΃f����6}�O��{�Fd����
g�S[���T�ƐX�6b�\`=f���C��sj�����ɬ7u��aWt1���x�8a�Ki��/F���j�_�Bh���{����'� ��NpU����UXWidi�Q2&}DILj��
?��K��<�	�^�{��i���1�R�>:�.��l�̇�T&*�e�̋ö�mR���˩ĩךS���Xe�����R��Q~�F��	z����W�ћ�f@��gRA�r%�����P2�����k��^tp���
uDK�X(�
)�;�s6��ܥm�6�%:!gw�p��8�h�#�IO<��Tdtϒk�َ�`��o�^r~~�/f_��y/�'O~���?���NS3GՔZ�[h�t��9ܜ��9���.j"SÇ=y{@=M��4�a�Agȳ]���2t��g�x�B��Oa�?�!�P�iN0��z�?��18,#1`99Xh��7����*,���L���:�mmRK��F��>����mGZfI���B�z5���sY吕uH�%I��vҀC\o�G���'xw|t�NTp�i����:h�w۹�����16Y��a�ud/�CP�g�fcs�2�福cz"^
@��܆���Ƽg�σwGT|�E��[e�Jv淅ex8�R8��U�kЛ&@\�S����|����ݺ&89�QXq�ߧ�܀4��!W�=S��h����X���[�y�e���C���Qy��c�?j�|2�]J���&)n�rM:|�H���ߝ9�ݔ���\O���8��x�"'%B��k5Y�R��p$�����Y�yO��8��Ot������2� 1�����	]?�V���n��ܽ���ge��"�(g���fH߯X`�u�mR.H��/��`�+n��.��v�lȌ�>:�����E�%6kL�z�F��ڀ����41��t����#������G|dF��?���SO�[�H;2P\�'E�ԽO���[��q�hA�\��6~�ì�#�,��*3�E�@���
J	��nҍğո�l����0�R�O�C)U�	�n�9v!e����-�a���L�_�]��PGJ��¼�)���!ϒ�.����*%�F��{Vf׬cm B,�ٕC~砫�FO����ҷic����o���uC��u^�Ȉ�h�3���HJV8���l�𤯹/�"cHo���8U�:a���9n����m/Z]>H���_�, 
U�\tC_�4Ml�<^��Ժɞ۵!�ufD킫.@jꓣ��gl9K�"mGx�����%�Y��()_�?H���^v^H��`�mG���:ߒ�?A.��$�����߰;��*ǝ��G��A���n�L���p9�i^&����=V'7o`���-��	�`�tRB�	>�ܿ��-��ä'm%��b.E�) w�����	k�C���_�4�����;X�9��'�Px��Tc:  ;����J����0�5�x�[�_�K¢}�5�r� ��/�}�};�� ׫���>��s�~�#c_#3"m?�K��Vu�-�`� ��kod����LkT�\p��U�g�W���f�D�iA2�=TN�,��V&�!�6�)�JGs#FXUG�܏�;`6$�'S�u���5�E8���~g��ɒvwɹ@�Å�d�r��~�����V�F�Z� �xM�6.���;�ƦJ�3��˱M�$΃��M$�Yo��.��pQn�7�!wt���+�\�xn5c�?�Wz���@�b�r H�����ieXϳ�h�FR�~X$��Mp�{[���K`�m=�v�s�ި��T��B�[.�3�xX�����L�b_{Lj����b>8;�{HUJ��
�8Z��/�i4�]����χMi����A�[̈��X'<���G�sT7���5z/FUZm�y�r.��Ż
�,����$F��T ���T�}^�T��&E��1����Ơ�6��bq1�ܣ'^�\���@��t��ZӠ�z1!��O�������f�;��	�ϋ���H�H/[sP��m:�}Kn��zݨb����� T�fAxXs�
b���q'ANX���L9���p�$�2����*m �����_[͎ ��/�6dmf���.��n1V`���^�ثЦ<�c����*3��%�9�;]JCK�RR)X<����F�\)�v|yOE@����P��%�(�<�FO���٨XlxVHYEB    fa00    1b30Q�4/۠nG<%� &?o�ڊU$�<#wL
��&���&#Ԭ��o�'n���A��#�<0�n�dx�"�]�|����B U.�~摠T�E�ʤ��5l��^�Σ��7�;E\�h�X�_/�T�Z��\pPC/*cb�����ޖy��J-5������D�w��<�"�'T���\V�e\��8D�Bc����6l��V�&9T���e:��ݍF�jH����]�嗸y���� �VU�}a*��a�N?�.��d<��Gr@�'��R9�F����O6�Q]�v�?��2�ڌ\x���٧�����yuB�k�P/j�|���$ش{˳."jy�_�]Cێi���//*�;�0�è��yz8O�|�4�,����-�`J��P�0@��"�_o:��J�Ԗ��:�4��cH�(�z����1.#{՚M������������j�/����Lza�( ��tԹ�N�Z)N�>�����X�W�,�,���o�"\��ut�E �X�?qTT��/�f���h�L^�9x���S���E�lMF+���^�B���ch=}��{�3f��a4 ��I�x��Wa�m\?/�c�49f��Q��c8�K�����Ii�[���Oɝ��z�Q�?���Q�b���������8_�����H��1���'��}p�"F�.�4&0���:�I*��p���>��)��B���l��Gij@�g��f��L=���G��Y�۠㾼M9������E��e*P���6�_/��	d��%D�z�Qz��I%����elv�vw�<Mc�:z1aL��K,�Xm�������T�i�6��Kg,�FGİT��(����]t�l�@X��(�w$���0��l-p(>Y�'�ܿ�r>{Z�J����(�$)�����v�S�޸C�ݣ�ƚM��j����;�h��]��i��⏇�/Fd<��eQ��t��@B�I�w]�\�����������0���R ���������[Cs9�,��`��U4�oE�aASU�7���i�I%��5���~���T�n�w���Ҕ�Kiݘ�T��1ܙ�k�D�eضh�+��C�s%&gZ��t�����K86�$rl����.s�	��@P�ݳ:	�6O���u(�w�	�m��
�Oe���1wY�^0婧�V�L���di.p@���Q�ۯ���".���y���zܔ�A.*ޖz4{3��-a������綃9�=:�R=ADq���uC�t���3C ��p咐�Q�����S�V�aQ!dQb���G?6� #���H��.�K���O-*$jZy�)�ࢤ��a�GY�u�i������KoŖkߘ)¥�T�����07D�-�ij��>� /ģ�2�ⷴ��JQ�����7���I0�F�%
�Z૑G~i�֩G����@$J����ЖQ��v�&��Ȕ/�Pրⲑ�دN�Jd�o�47����t��H+	錼�0�,]��*��ҩ�=���`S2hvU��C��ҔV@˵��ᚗ�밁�	Q�M�����f���*2		�w-������W|��� �����2.d���*1L��&0��ry�"���S;�r�g�b���l���5/��g1�`%�q"��t�ms�" T��*��,N�:|Nik��gg��GG���h$���B��W3n�e�����<T����X� D�*!����/� bC��2�r���a��*3�kj:k�n�K�@�m��n�	R���ð�Z� S#�5w����+��.`2��� �H�"�=�d�{^ d��y�/N��v�����`�"���{a��o!ʿ>N���m�¦@�Zm����2��܁i���69Ι|p����`'x
r;h#��=�S���f�Yb�	
8�����j����d`��?�X��h�PP��ۖ�;4וS����H����l�a*���]�!Ůr�BH�1$���b�W������D���)58:.��m<GW�E"��([?�:[�Fv��o�2��9��)��<��z^%XT��OQ;����5�D#|�6�� �
�	��ˡ���o=�ğf&h�J��<��负
����Hzs��}��yb�.y`��V�T�f,t7�O�&Q��-Z��=�Aw8��Ӱ��cf/����QAd~U
QM;?�V߯fG���W��G`�[�qpr� Ov�$�PP"7H����2Vz���U����  ӹ�H���S�
.�n��rQ�3
 ����v���:��� �M�E���a���n���� ���������Ls�IÎ
�������C��$ܮ�fZi+lmn�w�;�֘9����DS �C�F��I9����hm;�B��Ш$���䇻A��Hh��Ώ�s��}�~ވ����Χ�C��kk�{��%��F4=�?@t�^�뤏Gж>��ͧ-smْx��ר���z��z��_&m;7(�>�p���t�}�v���^��L0�eYƊ^��37J:+�l�,�oG��4v�1d`�c6	u�۰%c�;�gXh��CMh�O�F�h�[�k�F"O����f�S��� ��4��7�c���u�$֎h�P���?���c�9v,_5ϝ����~2�r��@ܠޱ�ã�<��%�ْ%��>��Xyt���fv��Ӧ�����F:l�	1z���G`���)L�7��5��
(��\+���3�c0��	U��U��OH~��Y&���Y�c��oX�B�j�v���/2��dBrK�Vj���k�cQԩ�缩a+���Ci#���Y�o���#���� �dggW��q�͛Z"�ˁEa�'�<��:����R��Aׁm*��.��f4{�V����1Ka���x݊�ڦ���D��C�`ޡ��ه�;!6%����U~h�T���ޚ��')��;�2�/�1�N-2��j�Q�𡩎b5Q3}�҄��$��u]FWI��as�c�_�KL쒚��|� ��t�є#��1W�<q�F+�i�C)@rܱ�G��0��>��%�Ux��-\�i�֧�\���L�b�ϝ$^j�����}���);�r��@���QA�����L�'f��'��fU��:�n�E�=�w��]΁C`]#�9O��Ձ�̣n�Z��N��;ua���)�3�R��ao`_0F���{�w��p�s7�&�;��$���]u�{��	����4L����z��Lg;E�s��|�c(6����z��6�˄�"�Z�[�&FV���`IF���w����&�cǰW�?�;�p�+��gf&.���$W���F����.*Y���
�eo1��x94bOU�L�C�i� �oD[��5�����J1��6[��X��4ƫ(W�eޠ+�l�<�>�?k������R*�4O�ƶ�߀�}� Ϧ�@`��alyݎ�����j9~��rd�,�#V��Y�P�y)7�}O�� Ck�{H&��=�n˜����ǉGX ��:����Y}�{��������c���Sx�U,Q�#u��s5�� �#�gyl\���I���s�82oQ���ò�)�,y��E�q!CG��V�����W���`9�6;����[Ǹ�W{-�
�/���_}�P^���6��D�`�91��sy����ހ��*��4�'�e�N�\�[R�-�a���iJz���p���頗�껻W{QE�_r�践�B��b��qSb:�VT�+*��Et�B���ԅ8l�����؝�)(/ݲ��P�l'#�l�ta�O���C��~ЀI�e��\{(9��WsX����~�g5z;X�)O�2S�m������3)�g$?%x�S��86��<�d�z���v�6<+5	Bl�s8s�
E��<[A@6�j6��Z�˳����[}PM��D$34Dx}�hTz�Rhƀ%5S��}�|�GY�ڒ��U<(P��G��^,��3�^2�ߑ��KX��W���}�r;T~�L�\�i&g�h�a�9�f�^��_=e0�c���>'+u(��L.���$��)��A�����<���~�MՏ4j[�K���(��A�ҀA����1�{ �eGץ��y_M|��9�K�=ѡәN�2B,ױ���wd��2�|��(�sө�If�吂�c�Ċ
�>��Y,��Z*����q� �S�a�A��~2�V����שe47i��pU���I2�#�qJqi��<υB>H���x�# )�yA'M�	������t��wx�:�w#V��t��eD^=I���%숈���b?�W��ڣmY�A��i�$0�ª�\����[;c��U[���4��a%�W���(7��4�Mڰ9ˢ����Џ��]��.��|b<�S&��2�LrJ应>�8��1��5�FPp+9���=w���O�A)ť���tL��T�Ht$ �?iؐnʻ�3Xhu��/ɓ��v:�r���%�x�{V��0��f��4��BI�P��gWq��8�v�s���ڔ�on�s�����t��(pO!
�X3C0�!!���$}�c�� : x_�o�Ycٙ��������{eXj���ޟ��
��b 1�>2��RV�J��TR�����|6��1�٦�&WpLƣT#,��蟄7m���~F9J�
,qV�q2�Z���,L��G�9:��B�%̍�Nu�}qN����������m�Zf�%�U'd�w�H���T0K�űo�g]��vT�4�d��z&�ó���*��U̧���%s}�8\Ղdd�B�6	Q�d���ը{C�M�ۺʵL9��2��=�Z˼6Q�Q�0b��@�3�0@I����#�Zhѳ�B�;/"u����p�g����0:��2�GkͲ�_���Sn�~�K9��v>���j��e��x�G�����^�!�ũw���>�1��\�����f|@H `�4n�4�c�����Aܒ
��Ŀ,D �%��76�4��\|�涫�%o��A͜i�tVV��]��X���D���6ߘ7LXD�3�E��l�$�>���H:Ey0͝� rYVu�iM�����p\��9_�	!Os�t���|��E�k��4��WL(�;�3_M_3�=��%�*���p0�����v>ش�rOOL2	]�G�K��'3S=����c�Na������٧�꼿��7L�[2��7��/�Xk|�_�̸��LI�x����s"z�תɮ �Kb(o-!�c�d��Sf#�`�6�Z�_��1�tS�%���'Z70�S&�R�-Q�o�F 2�1�oR>���;�����vr����Ҷ4CAm:��+�~Y�Gd�? ��u��+�eT������|�bX���S�yE����,����|��G������;l����Q��ѝ�K����t �@c�#�gd,�NL�;��9�q�>R_�wᓅhX��~�]�$�9�KokB92�0ߏL�C1�a�}*=C�u:�&��=��\G=���nHii����N�M���.�/O�g~�W��씷�c~�<S���)ט잜{?:s,?�Z����#����� 7�^�E ��"����Pczf*2=��/��N���Yy�V�'�� �}�?�����.�dIG ��~x�I��Jr�6h�8Wq�8�Bt��֮�H�L�<B#@3��CL:�<�#�:������y����A���4ԃ�G>��%x�Z�������5��V,=]T��G���d2�!�Jg	� �(��.�A�)���w��ē]�zQPNA�A�z,]��ODIp�ȓv��4�8��0*@� 7��X�"��ȅ��
��Y1}0QJy"�_�����ꐗB�4�*�%�C�Ȣ�IY503������=�X���%�I�`Nn1=�2�z���i��m7/�l���ҿ�Ă[ۦb"kK�p]Hva/�'U#+��zP$��>�$����Z��r�#��Սy`�O ��.��E��P2��~>�e6Q�v4_6GOQ= �A��o�N �"��[<��s`�AoN�!3Y/��C��>���=��!���5`I�@�?����'���jt���%pSt�ίC�XM�K����:ob��1x�qG/�Z��� ����Ȁ�u���r7�VgE�~�5���ٌ��v�vG��\�0Jm"�*�[;�B#���;�D��y*�Bc�-��?�u5�A2=2S+V��/�4��	�wD��O�r%*���J�
�oM�u-��r�� � �ͥ�?2��_~/: f<E��"���S	_Ȁ	y���}a^�,��Ȑ�+����Z��_� i�Bzm�_��ׯ��3-�Q@��?"�=�5|]�[�D�L�ɤS�%�o�� �feϴ�f�m�wޱ5s�������'EN�j�/ƦP6����cc�*w�K��1�o��A+�:d\g�"�ˎRm��G=��j�U
���HМέ�a��rSU6w�=���!�9�>���u\�$\B�T1�T]u{"`�0������]6X��.��j��q0�fw��^
�ZZ_�B)t�����I
!3-Y��V���Mj�C�N�u[���*$�*�( <��jߥ���.��h�ؔa�� ��q,jʵ�ǅ����˴��K�`���<E��6,C�-K(�j�\��X�/|u'`�]��I&,ֽ���!y�����f2�$����(�-�@�q��B�2�ϚD0��}>2�x
:�1���N����%�<ҝQ��ݾH20��~k��u-l�L�Z�$ac��-���W�qV���K��8��b#�7R�W�n��S�D
�E�X�0�wQ�|e�,��ީ���2�^��j�C����[:`/8 c�L���(vQ�A+0���K��X"Cf��iP�̚5+��b¯��
[����5 Mƴ)�e��θ�$�R��!�8_-�;�����m����XlxVHYEB    fa00    1950�N�=�O	���'���
a�������β!%k��w������9B��&��@H����s��3��A�YD�'��,���%���T�*0�������-���B�H��r�5P�-!���
n��!V�&Z�1�����?\HKUs6`b���n�ZW���&D�E*Ŵ��-�(���-��@��@/3/�=�Nk�E�V<d19�iυU�?Z�H��@�hM�l�`�Ո��ɼ
sK�ۂ�4� Ma���}��Od�=��R�*%���2pU��ώa�}��ۧ��͙u�k���b�3�K�j=�eVy� �p����v��"q�L��3����A�l����D8����9ߦ�t��f��cCh^({�B>�K�72��׷�
f�a���3��Q!w��	9仉��P^�d�r��%;�W�q4�VE7����E��ok�s�h_�}�6V'��g�U_���WY��ŷEpj�j.�G�V�ڻ��q�]�t�ܲ��@p�9	�$?
h�P��WdP��T��<~y���qO��1t[���e�2����J]}X�UU�"%G�9������n�Bݝw[�=���UP���v�v����W,F��G>�\Ӓ� ugm��ݮ���M����O��~����?�$�t�W�S/yK�v�g ����L���g�FC��O����I��3�`�/��J]�����
:�	��jƷ�Z7�	�F���@�(j��Q����kw����,��N��@z��p$��>ơ$\�>j1����B&���E�;��r+�N�B�A�:�)�|�F\,�W���@%|P N�r��I�3؟�6$9K�|�f,�Z| e 1/G�%?�=d�"_P�zW�Z��G�O� �x�F��|s}we&�
��Ja��_[�J`H�>��=���������N�=?��/hm.�̠`��"c`�T����\��x5Y��۾�����g�H qvs�wp���غ�\]�N�^�@+�Hϱ�	��=�a��ڼd�5W:ja�C������Z����{@���ߠ�t��"�}{�$|mѠ:6���:TrG��r?��K*m��l����b�.2@��2�]�/i��}��t��7��z�Dg����p�7�lmM�����/��LD3}T�}�	6f� �N���ܤ�&'�VOt��2ٳ����Q�C,������M�+\�~�03%X������2�̨0�g�X�����i5�����3��.Z��t]��N[�l�A�Π���z�,~���^�:�8�/q'�R�\K1V�,e�r!>��;�Ϣu��Z(R^s0�=d ��(k���t4�z3��P��l�$�
I���U�L/3-Du'} �����Rp�?��"5/�����q�h!�Pu�;�g�_�.�=w�#��<p��B��6<����'����WI��G����;�\�P��3d�)|���ݜ@O{V@M�\��Pe�+�W�K.�	���&��=85zu��x��_k7��%����2
���D�Hqq	�r\�y�s�����s@p��Y�1M�% @:*��T�Y���Q/����ǹ��eFn��Xߞ�CǨ�G*��22�-|۟� ��7!���*�����ڋ��ll�tjZ
����[�)sˎ�����G�emH�L/xX�Ȝ��_ָUT!1�r1f5I�1è&.ӌ���*�Rb��O�7sθ�JW�$M� j ��IE9��ؽӳ��/�脸\�i��l���%a��`r����T���/<��7�Z�b�1��}|%���(í�f�|T�/�	� �:M�V���f���)�g*]���M�}��z$nüa7N'��C?�W@Ѵ�tV|�F�\�'��#SU6��[�ʵ@�� ��?j�C�p�T���������r"=�9����b�`�Y��ivNz��C�FJS�&�0�nTM�-�~��2�d�|b���9��������p��H%/�ȔtJ[��*��Ι*\����7�
���mkTe���)�Vu�/��̘�[�0X,-B��
ש�j�Hy�)"x~�?���&��{[K������f
��rD�&��^3i�X��m��
h��`*��ԿWDWn�É����4!d�PUHEwN��I��AKN��I����q!����3�d;��!�d�*�T.�s�>�UVq�瀒&拘N�&TҜG�>C�X��?�1,ԑ(����)o��E�[3N(�&E"�~֚�����h��)�����;I�e��6��+8�1P$n ��9_A�k��� ��"G��!M-�O��*V5Α�dt^O���N����@o�ؓX��i*m$�F���/��Ř�J��Q=��}N8�N����'k�J�s���k`��r1����b��>�������J�/(��Q�h�js��cSu�O�����k�"����+굝���U�5Dg<���]��<:ʤ��'l�	C�?vN�,?|C]��{��)��5���	^���B��`�;�6�X*��t��p�$5�h��wS8��X�0�l�p�o�4�% ɳ���C��[ ��(�f���ްZ���+*�؎��r
��:M�8�h����?)[4ǜ1��@�s�zS�?�1;+�E���f�>Ĥ��� �6x-I�NN�>�Q��j�ψ�8����z^>��hbqRf��蹿�gW��n�-9�D$K`yٌ&(�����
�[=t�P�Е�/Ϻ|;|��q�d4�4�R�P��8�(4/EhA�օo���� wN��h���jH��y����md_	juYl�hb!sG!�_`��]����n?�E�$뽘�w�p��0���*��� �㯴'Po�#���UM����4꒵�?S��$0-[Ui�-uw5yOL~��% R��h�M��V�+m��j�Q䓧���<�#U����|K�h7��w��)L�~Ea|��r�'����.��9b ��.�1��e�1:�E��#z\�+fN엜��b!NA��s���/6pXh�BGz����e��)����`Czj�)�ty��@E��z�Q *����]Nv��L�8+�|`���������!��a+����p����h�b��(�g���.#V�Oz���(V����)� <�.�<iԩ1�s�
����r�U�rFִn�Vd=�L�81��iu����y�zH�'d [W�.7�U��)!�p�ꏩ�%���8.5�G�h���,+Ϛ��3����H;����V~�o9d��Q�q#=��`�Z�i�yK:8
�:����&Y)K /|�'C�T�Z��#�:�lw}�h��|*��Ȉe_����zΔY�{�tA_U�c��K��	���$�YHjeɠi�.~E8�M��gxH~�˘�ȺU,�ʌ�w#��"K�5I��␜\��Qstd��)=ݸ5��y�x��R�?L7�1��3��/c�z�;h�^3T�s�e���sdj��1������D��C�D;eX�qU��[�����~�ƫ1@�МN�0��Yb.��v_]54h���S���4�>���'ҦD#�iC��m�?�=��4��w�3\"}��᭩�����ּ�3@�s�0������pV��96�@�J����|3�,��o�ø��|�$=S��+����R��BK3V�;q�O��9�����=�I��Edytv�o��T=�sCL�-�`�"�F�NWeb���o�
�~0�=�x�9� ��S~����NYL�1����p��+%����W4�A\��⦑�� ,Ⱦ�������z|0�F����P��\��C��C�bHP���{��*�	n5~�< ����y�[���d��(�z��[uI�"(Ȕ@��n�)(F:�Q��Y��I�恏�={���}���?f�;�c�I~ 6[�4�;B�BpP�N�C�kR�J�ZURj�����b�@
���Af��dI�E�x��J����	@��C�ɞ����#Z�(���,,`��۬]���� 1v�$��%�CeN&¥���$ya��I��	d}3�����2Α���^h�v��:S++80ZĮ^-������}}2%"s��D�D~�E�[a�=a�t[��{��Wr��ȼ��F�/_H�����J}W?q�`G�H��m(�֮��e�P��:C�3�6���!�����+f�ݝ]z�[�0ѧ�H�7A�|���..��Iy�D@��N:�iE�}z	��2�>����l�Ԙ|����"[]^q�|3-��6��5΀���~��6�W.��?��"�X�P�^f�L&�Bj���j���"?K�I>3�%⇌*lw���;�l�UOH�h:�̇ ��e��y���S�c�%���f�3�R�ӑ��9�![cG��I8,�X&��W�PNA)DȌy��8��P.#�+� 1 '��'�g�ڜ1�u!�:լ�0��Hi "�~�b�$����@D���CK��׆E��7��Ж#A�u�q�KW�����I����@�b�>��6�KEtPC"UT��������X�q-���B�]1��f�N��*�)��1���!� d��6�!��2�r>��Ɣk���,$��V3��Ox[�����Ke2��Zu�R���*��qEo&4o)���P\���8��Q�I�E���x��CV$�>\��b-�w���B_ʁ����ϻ �K�f���Mp<�`X����+��'��}�[���t�Q�56<F���'Į��roɄ	_�<��̿(x¶)>
���iO�:ө�%;.���`פ���ޥ���6N2�����} ���*��&n�X��&��(=ٚs�#��ZȻ�-L�ȃ��ް��	�<�X�^����eX���R� 㛕x��R 5y0Ẁ��8��Ɋ�aU��&eW�?G�8�c��h��� h���*�Ty~G�m~,�|�/vZ�\������M�g�u�[��>;�0T�ݴ�"U.�g����F-����=2I�Y�Z��C+��	)/�-7���B�5����̰���kI�z��o��M�n����2�����  -Gy6=�T��T���#��,;���6�[J����̓뤝>�\���{C��%n̝��ùYH��g�׿�����WB8tg*������6<���K�acn�hƥ�j^J,wo���F� �"2��K_�h���������V��x����#��{�?�S��N�3�X�����Џn[�''�M��9I�q��~���e��7XuG�%��~�.��mc,�YY���d�*3�omߪq��KW��(�uGs���Z	���Q�%=�l<��%T��||�q�FL���~=��-��UA ���5�����Pé��F����& zp�\X^_,��r' ����~�
�%���Os^m�v~�xL���ҷ�����,����B����I��H���xl4�6�-��ېpڅ���}�$B�4m6�e.�Ϻ����jO�	��:/w��4Q��A<r:�9����"��Un���y�w'ިNF�	`7��Uqܟ9�G38��J��>�>;�|\и�&1�![��^.-\��k6q{7-��5�hq�a-��	k0�dV�م� ��Z*���t�;�|q6p{(�]��TC����p0�_��y�3�d��'�}�WY�U_�v4	��;����J�����PJ�(���v���>߻���-^b�sT��V�Z 0���d.z�x�eg�=��utHYV���dfo&�G�f� A�Β
��߱�[��~h���N�� n��Pg�Q8�hXW(?�a ���k�b���7gf�5��WīƢ`E�K]zm5*d�p<�9髣\����'"ܬ��=�$���p,%�b9/Y��`�+M�kٰ}�+h��A�
F�����⁠�R =TRϱ]���=���Yh��lTJʭ��OK�ڠ�qC�Ż���׆�2V���}����H��Շo��ԛ,y��M���]�5_����/�Ub�ӝ��N�k��� �8(c5���6�6�&�wm5J��ce����e�hh�@f�֋�/�\+1�l�[�xV�������%(t\z �K�s4\���T�g��p컘���!�4��2$��A�Z,��V-�d��t=�]�Qǜ�
5O��r.���%{C�O�Y���Vnp5���F.�y|I�B�[y��uGm�����#���g��3��]R����K�e������D�w7���6����X��
�=F���+�n�	N2z�woFɮ���ԛ��1-�զT��^�)T���T�B��R,<�B&�5޼NXk15$�Is���Q ��#F���T���PG�Õ����=�M�f��0b��}>;�Xn��@�{Q��^\XlxVHYEB    4f27     d40198�۸)��}����Sp���\]֍�3�fP��v�����:��/�RX  HP�k�/,VG ?����\���Ĩф��d�W
�Yٷ嫷=k�M����=xLZ���u��U����%`�w��]wL�/_?bډ��;�_�a_���p9� �� b@�Y�d�kCZ������q�X�$Sι(�ˡ1�
n�7��~�~�m��*��=�x�ֱb�*K��V� �X�H C��v�j��&�t�n�ڒzu&GO���a��УP<��kp���z�N�<�ֱ5�R��jQ#8{�E��WR(<7?�1�Y4��+��^��8���M�'#�bo�n��Syw1诗r���6�d�nlB?��Bx[�Eqg�G��o���ʺd J����,���}_��Fn�+�Fp@Y�G�o�1s�^�I(=�Ng#_�\��<�oc�?c���^D
�]�̲��'f�}���7��6��$X�0����KѶ�e�E�F�����F ѽc��MC����!#�P w����6��-�R}8Ƕy S��	9�FCiMCV�|��nZ9�|���$���1�Z�u�ݝ��+3盎�S���z6A��P�	��;�:���㴔�R���M�=����5���s���Ip&��HK.�N��'��y�T�,��}j�k��R��+�ʞ��rK�����-�,{�&n������8a󙿠�r���~��<�@ڥuC ������,�+�>������[��AL�,�V|ԡ��<.��c��0�8 �e�6�rEw�������gE��0��uՌ��W{�vio���"�+{{�ַCCY���ok�h߂v�q��r+�)4>Ѣt�ץ�Ԗ�(�X��p��e������w��Y�=���*�N��p��P���n(�${����,Ke����R�R�c��B�Yo�0?<���k܈�e�O��%I����\Yn��^�V5���=f���	:Q�uHå�-p�[]��T����,C\���݅P���u��E�K��Q��$Z��Y(�mĿ`eL���=���hV�-ｏ�܊����7&^4�-�#ٌqM#A��E3�fs��:)��5�������_�ezdmv�H����<8�~I�Q�KCHn�\���!l�?�˶�p���8�� t0����57���y�*�����Wﲄ�[r���vG�t<��O�WR߷Ӕ�3w�cNC�Mo5���&�]�6�}�bw�-�>H"���E�j�=F�����Y;�'��k��t��U�v��^?L�%��BuJ�I-����l��rd�#2�f�!0��;�Wr�k��_���@��ҙLuX�B~o���2�l�����&�Ţ�w�oo<)�jV���z�n2�<���|p�z� �������z�<��)2��Hl���ڰ�`W�h�h�첯m�]��18f���v��/�
84'���T�w�U}M(�qcL��\˒��b�N{�FMz����kZ�Z�G��'����`N�d�K/��wU2K�cI?����Z���N܌��مb���:�i��Li�#O�Br��j�_��ޝX!�>d]c2먃]!����?,xA��6�ݣ�ώ���������(�H�/��H�.%S���5'��D�e���*gQ�®s%�#E����kΩ8��V�n���1��!&~#�b����E���Y,��T[�
���>e�e�&�-F��6f��m������9� ������rZDX��r��u��*��~�����&S��a�Y�h��Dᘤ�ߔ	D*�ce�s��U����$�䖢<V�h���Hft�dꈆ�*��Ѿ���H�ʉ[G��:�A�SzA����x��������QF��p��Ґ[5�.��8oUMEZ�+=a<Uf�V�:�%u@Gڡ���@�f�5I��^M��ƌG���V�Ƭ?o}����YAQ}�ˤA27��������9�+�x���?��טU�b@���
ί��T֧x���;T�`q��
\���>��Z-��u(�d�����u��X��ew�L�e��Q��_U�r���@brD��J�*J�$8�a\_ɏV���ў�I*.ww�ލ���^S�h���?qҠ���#��մ�?�V��BY:��.�D��c��J+��n\�N��	7���=Ӣ u�:�M8����k���q�s(Ӄ~����M��=[�y�|x��W��t�.��b�^����'K@�Ҍ���)���|WN Am��D�*1�7Sq����t��Dѱ�	(CE���mU���`1~R��0�O��,�L���]��^��=�/d]y�I&�\t�`�	=�=������Y��_!���&.�a0���%�v� ��ݩ�20�3i��&]q"�����z��g�P�#+�U���Q>�:>�,�\2*u��Yn�����2�7~��_�rs��������85�R��%Q�T�Y����O�S^D�r�O��E3���~"�kt>���F�t�[��{N�iu``��vN���P\$�1n�L��Iy���8'|�m�ˈƊ��y�T=!�.L4\f�ú��O��Y�cw�O�C�z*�~?� ���
\�����N��C���s��Hе�:cu��(�b�Z�e���y��uO�+T��?�������(b�ty�}��ę�D8ȇ��c[%�b��[EB0������p���c����� 5�,N�1�r��ԣz�<[M8��Kx�U|@��9�Bw���u�&�QYd��A�0��a��[��줗V6z��\��꫌1�s:>��: |Q���O�f�6�>���
\�8��Z�~}�E�xd`�����*�
w��Jr1�����aֺ��3'Pw\2�1~�e$|�2�����2lf⿪��<�w$�v0h�{5L;W��[	�P殻��gkX��ٱ����S��@D�l��C���[�7w�!�B�Gr�ٙd����Ti���z�%�:\B��7��!EI�h�����(���gʵOs���>�-3�R�/ ml�dLC.�_�z���o/FX�ȫ��^{'�"ŗ�zYP�]_��k=�@��*���'�!C��� ���(+Q�N��r���!�#��>w�v�Ѡ��_�ئ��V0K��G]���Se؍��}%�A�� �����Eޠ�~zz2�)�rRT�ñBvb b��CK��]j�}��oJ���\�S���_
���9i(�ŋ�� K��&4�Wa5߱RJ��w�ޣ;S:������w�D&�dC��}�-������t��E�E�$$ŎTL�a�;dև�ǻ�Zai�f�w�c�Df-�U�`1� o��}���+,��-�"%�