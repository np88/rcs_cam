XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��L�F5����95��~�~B�H�z��ρԇ��}���x�?��{4����-L�$ߦ�� ��|�Q�ȋ`�񴣃�sᬪHLE�$H��rŉ:.J�4š/�"��� y�F�Мa�
�T�2ʭ `u�m�="8�oRo
〱Q�m,^��H�:�C��t�i��V��AT��K��	۸&�蟭�����@�-/޻.�Xm���H����Uk�+����լ�J�0~�C���&�a�q�sz��}g����0O(y�ƔC���åM��^�/`��u�B��zSӗ��D�a��`�Qg�%ٹ����9<ne�>����oJm��bO�e�F|����ȯ�� �-���&/cd`��×ȏ�hM��ILA=b"��՜���������d�+xQ���n&.�'!Qa:>�Ŝz,��N>�(��g!E^ܧ��D>�`���j�,�r$ڒ~�2 ��ȌvJ���h�2ȶ��3$�&%5�����6�f��<*�E�9�Z��@|b��y�!CGq#N�J>�3���mI�� i��,�X�z���']?!����LN:�32��'�E�qя.@)ʓ��y�[�_�����%:>�F�
0�KUZ�>9�Ʒ�Bl{u�n�ݘy�$rs^��a
�f�t��H�q��Q$�/�i��H���~-ec�~�W�h�F7���a�,X b4�?N����|Ȓ���<&���a�1�E����α[���{PD丛C�9]e�kx��@�d���ʹ���Ќ� ��N�&��Q���.XlxVHYEB    9732    14d0���(5���(	�̧��n՞fd2J�����8a_�p4*Ǡ�_��ލ78۞y�>�F��n�����I8�l��<5�
�8����ﴆR�����U<ye�[n�X�r��~Ҝ`����U�. �ⴵ�|��;�2�D�!'+���\SX%cD�T&�=�.N'γ���*Q���w�6��æ�n���T�/��gP4�}�1hd� 'y��Nj���ϖJ��cm����`񢮧Q�8F���u�e���9������?�pHe��N���{__��[��M'Ŏ�A���Z�� b_)ſ�uP��Y�P���Ix��֑~��R�x]SJVH��9.���1�J����,�!��f���ˬ*��Ew���؃�
���rz-ȱ�廯c.&:Z`ie����t�%뷭�r��%�36N�3�t>?�3�Q�O}A��,���U��Ye9�|%��<���ޱ���JC��j�
��6~/�;����@L�2v�3~���̐��m��������=w-��l�L��3˘� �����Sp��6N#�Y4г���ۘ��&<�=��꽰����2����5s�F;6����D=��)q��LPR�p&PI���c�r�>��9[,4�-*=�M����?��R�I�_ߺ~���&�ث���j�y�RF�<�Y�8��z�)���+'�J��wZr�������p�]���6OF��Fܜ/���N�]�>��5k|	�`�`��#:`J�I7k�7��z�v�-Dhj*E�L���m[V�Ͼέ�ͥћ�����ս�'�PCg�R�U}���?�4��⎫qp���t���JI��Z�tOnJ:,��UI���q��8���	�mQ�0~�+~ħ�)�Ђ^N��<�ͪ���D��Zn;G�A2��Z�A\&]��j�)%sW� �Q�s��y����@��[�>�Wui]-��\6�%���y��ӓ�J[l(R����˕�K)�	sG�s����G�cǾ#�wi��������r{���hC� �|��Ҁb�����<�z>�FxL+�763/@ھ��j��_�e�|w�|��)�%7ڨ&�7�
D9C��m�4z��`G�UB�o8P��
�[>�����~���)bgT;,A��}ir��p�|s�u���xW��4!b��i^����RDαk�J��:S�P!~gu*������?����)p�N����쯑g�Aڒ�9<�6$Jj��.�|p�5��X,ȕ�a	�wz`5�Ac��vW�enQ��K�]��c5�70X`Wt�6M��"��Ӳ'��j�4����N��������(���W���W������|-�Q
���b�MZ%zs��5��f����ń4���}>��i��p��7^���� |�����LY�"z��{=Am������yZ@���j�̢]�F�����:��<� �/6N���*�e�����ޚRT��dpl#gYN+�w�U��6��Q�%TЖ�?�[��͟���D��j5�PZ��W�n�0������se/d�|F�A�K
؛� ���tSJ9�\���W�g�ɧ�P�(��/�B�Ϲ$׶h�P{�/�gM����w��5�w|�۞5.�]"���Jz2�F ��jZ�܋��,�S�B�̝���y��1|�-�E���i�S
��}:[%�68WlO֚F�v��7�ji���?D]�Y�[���+�9��@�����Rf��� ���_�,�i	<����W��-n'P���:�r��>�C_��zv�cT���(���)6�oP�����������Qc��ݬ�?*�x���d�^��#$����Lq�Cs�ǌ�3w�@Ѫ!l��Tq!C���E9��}"�;��1��r�ts%?������.�_���iY_������Af���'	O�[�쑴����k���`�`7Y�(�:��:�S]�+��W�l�ܖu� ��F���YL�;! Xτc���3���y��<;��L��T|���G�6��k�]���w�H	�c���t9��\���R�h�)Nb��]��B� �����D�:[�hƾ��
N�ZX�U�"ظ�\xȴ~�O��W (�8���������� �C�_���<����B�f}�s��L�[+ɲ(��a�k���+�m�5�9�,
1#��#HH4��B2�1�Q"o(�ʓ�`גS�YXG�����H0��^n���[�::إ\�H؉W�����m�	����s�f���?��5v��cru%1��Ty]0�T@���m��0&u�����1�W�i-5��Ux���:�����yYg$ O�>r�"�����A&K���g�&�/@z�"!��j���:yb!��A��J	.�.u��OwRZCP�=�DZQ�"��N�͋���y?�չ�'��o���w�sKQ��+^��.��@��'a�8��)�};R ܐJ�-���Zp�k���'c�ؚEKr�����
i6�I�xꇊko/������>ےE�R�V�Iu�U�K&�!7
��g�MUA�^��h��w{����F�-A<�Ĉ�h�+�]��)x���&u�T��@��K���I��ut��4� �=��[��"�A��۹>|���R�͚;n��%�g
���_�dZ����F�zr2� �e�s;8ˎa��pxMD[�U����[K�h]�K�Q��O1ۙ����w�|���kp4���<�"�h(�
���#�6�	>L�Q�ԛ�r���9i�ˉ̓_^�ct�clA�i�zh���e�r5��CT�Uќr"^*����_ckw���7��T�ěbZ׵�
,��]+�=Y����v�V���ȕe���e�?$ߢ5�rײժ|�]�I��?��i"�'[�f��' QC3���Ǜ�+��B+C^nȀjy��D�*�I+77g�3���4�f}mn��\s��7L]r_�"�u��_��׎0 �4��]-"�7����	�d�~ʐ��W����z�GZ���3\���.yl��7K:���0��̴�J�]c9��z��2�?��C�����/����x%7�c$ٵ$��A$���/��$����~Y���NZQU��Qi���zI��~X�W����{���J�md�o�lg������nYy��$wտ��T(a ���NAr!��O��j)F&����L;��Ex�b��ⲟ��3
ʹ1�,8�C)��A%+��v��N��Ȑ�_��dZ�?�V)N�!�R�;��&X󚭚l�o)y�i��ThMD��o��ML��D�hY�E�g}���-/�S�-`���\����%��J����}�
��ϱS+�ԝtì��S�����	K��� �����'
�c@?��b�)�x�c�_��T�X� `1E����^��2�x���Ie�T#��@��{@�v���j#7M�|�y��=��S��x��p����t������o�U�^�	O{6s�4kĩ/Ri�������)�"�8kȇfNx}r����i���\�� ���@���0e�7Cg�i�u{���m6J����q|����\�'�ݟ��%�r���-���)t�O���)�-��"t�cA/]?�_�L�A]ja���O�X�M�o̜(4�xK+s��Į��U.֜ZE"��>���wh��!'?�W�=?�J>t��^��f��]sʶ�K=򳪳tU�j��7*�}<j`���2<��S~��hks]J>�wm8J20��e�c�#O$��?NY�ʱ�$���ߵ~���ו@K�B�q��G ��L��{�̈c�L�ii.��X,����j�42���0w�W.��@G=�EnK�iA�:i&�
@ 0ka]3��?П+�G!<�t��Rs̹ ��6ʥ,���8�s��FWh�uE.F0�*+X#���RR1J�����Һ�7#��x�L�HBt����(�/�񃋟pBBG�Ւk�
�9@`�I3(�[��1�.������71"��T���;a"([���=u;�|������bدX�V�u���I�7���4�^�#���pI'�E`սοS(u��&1���������ox0�jD'3�{�\G춞g(�*�Lp�n�g�w�Ew���nn��S��9%^���������5��\0f��������Yu�b�g�I��uj��Q�0c��z#�	m
��
��Bf֏�9l^�$���(k[iI�t�����E��%���'���A/�{�^@�.�1sq[x}1Ǖ�e��X��¿	���X� ��k��yQ�syѨ��
%�y�&Í��7.P��s���8�c�mf�aV�M�uA��%o��J�c�����sK�+D�}�,���궮���=-T*pu-e�V�i~hb����5S�m2�����jנ�"Ψs8�q~�q�=x��ARC��Rb!o�^D��>��`��F��܁�?�����Q��b�3wV�= =q����>%�H����
����H�2pg2W4n4�ͯ�!�4Erd�^8F3�k
�!����72���A?�I�»�)Iɧ��ӥr���x{�)��V�b�Vd[��e� �I̜����K=�޵��ev��7Fb�r�/���
$έ���n�#|	 ����r9���p]!`��DեWMԜ�������FУ����+���&~:�C�ꑎ�I��L��9[��pI&|�X��{aD��iT��^�D� �W�Wy}�[��R��G��P��:ޫ���vD`�5�<a���9�Lnz��qz��>�,�z�[�~�%��)��#���	腿�sŪ��O#9d0x��+}��۩C��_y�[��%�z{֪E�0p3@�v��CJ��f�	�Q��A�X�<v�0���;�t���c�� ��s���gM�Of� � ��[0��b����=l5/N�ɕUz��X��t�(8�bJ��t��)�������a�9_/���g���U�U��xŞ���{|����t>�B�,�Z���,�C�꺦/����_5��R,�jet��R0�uТB��&^m�����X�Y���O�!E>i��4T�+]�>^օ8�$L�k[f���J603�!O@�OE)5�7�K`d~!�~���`�'IE7_A���H��3��?$���gy��љ������f&z�n֕ �x�xGm7R�č�6R��Eh{�3A���^n��Cǘ3U��U��nw9B� '�~+�n_�a�C��X��	YrH��軯��L0��fp3w�4n�OQ��ԡX� lv������nL`b