XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��k=� 	�8��VqWI_�����q��چq�i����g��J=��΢rn�S���ʓ-�)�B��k�#41u��n����>�A��3�s2;t�������Zçӊ?����ĕt��\��X{Ʀ�rw�2���T6�̙�-:h��e+ٜ:��v�xc�樧n�T����RT�GE	
CD�j��/�P����f_u[�up�ik�K��I�E����榧Q�,�_��m��9��6��禎tH����8���k��,
&�-��4W~�}�1S)���]جaa�01�v��TA�j3�Y;W�V�j��������U֛����*�;��g]V^lA��b'h�.�n�N&$n�v����b�U2��"�G0߀Z����˫��q.��"8p�Y��3���i)tb����|(���WC�b���yհ�H%?����9}�����'����K���� *qc��m��.zmU�ۭ�|��t1@���M�El&�&1�����ЃxVE�fp��ǃ����5E�)}�	&U?�0�rCB@��	�cuf̫<��p�X�~ B�2p���������{���zvx�\��E�7�ݸB�z"��+L(����b�q���m_����"�	��(��8���,Gi����:��1�IT4|��A�˄:��}�h��w⟘�t�$�*�a��$';֡4���C�>Z�Hcm_8�����ݎbf[�O��b{f�D��ή*�)F��H�>� q*�E XlxVHYEB    160d     7d0�n�,�-O��}�_3��/9�QL�,]����)��K�͍��/�76��� ��V7�W�ĥf�G���S����x�G�����C��R0�
� ̣��j?�4�)9�wqus�a�Bz=��$��
�����.>���@�ZY�#�`A����M����:�Uj%*� N���/�z�	��I?�'z�q,�5����j>[����N�>��zn�W�ǂ�7�N�4�ї�QIlQ��|���aJr�����pz�A�WQغ��hp���Bp��)Wd"=�$�����Ħ<�NgKQ�&Πp<=�G�:��wBż�w{�z�#'�G����W�{~:�߮M�0c�A;�+��j�;	��)�:�Ug{6����H95�zWU��}n��(�WPA>��jW�)t�0�؎�ZE��݇���
��U�P��x�k�3C$^sjHV
(;�դ��[;G̬u1#!ɪ�a$�Ӿ�')0��J�*�R ��!߻���b^h�9���3̹7N��l6��	l%���{�R�~+�&�as��1�v������3�6������Lf������Ã���, �չ�s�x����z1�rfA%�I�/�jI	���pV�_;�(�� �-��I��|+m��C�զ<B�~�.'����-���1˂���S�l%k[9��}���&�K1�aQQ�k�0�K9��HҺ�X��Z�"|"Hf\��#�hk�_C�{R���&��4B�.�������^~�ݺ}�Oiy����*�>���.Wp��y��ూ#
��7M��U�%�߃NT����xc'6�=� ��l����}�T���y=�*�	.T	�!>�Ym�uA�]���i���0D��mi��|�=V���a��G�w%�@9�Je��=1 ��ȯހk���̜��5R�
��*H�TS܂o���m��q,u�;)��uD@p�,9����8�=p$T|إ��T�RĐr�U~�����<������O�o��]Bk O��ġ�H��h0��������UܗC�#�%ɤ@m-�G%��L�~�GL�ȅ�a���T�w/*D\}������;<ƶ�~po���Z0�za�a��w!`{g|C�H�}�o�:h2���\��گ�5d�M����B����2��n�[_g�hY&�D�N!�s�/(p:���N.J��ZX'�c�'�U�o	\�;����]���:z�"Q�/a������~[�Cw�3T�;�<������eFͪ����mn,�z��O�DEt�k���#)�􆴒!	�����/T�C���W=9��?@��R$^��Դ�ٖ��U�e���PY��hV�x��T%�h %���Z?��Ɓ̼�áD=������p¥�1bq����	KO�&��lx�Dą1ā-��6 ��\v2�a�Bs�r�NO뎲��!XH��*]@�d
h��[�x�&��WBk��w�>Ae��ٱ�t�Or��Kݳ���j�X�ss��}��O��,v�*���7�)�VwՆ�\ږ�X��G���MOO3�6�gG>��#q��z}�c�����*��_�^��=�]�:�x�yKN��BB��1�حԂ; �\�]$ia3){�]���T�TnK��~��e3\Dw��������s��y��P��f��T�Y���F͋��h��t�>P�J�.*H8��	�O�־�z��)[��0�lQ�}���K4��$v>]�Sʾ32���>iݛ"��
���5��V5#�Ȝ��M|�]>䖻���l�Q30��� �o���z�h�e����ڈ���'&O"s ������lC')TG�*�Ze>�Y$(W34�R���ߊ���쟄@����z��?;���!���8�w�����Hob	��݀FI������
�ޓ�ܪ�N�~W�F0��XlI�B�0҆��,'