XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��R>T��m�<��Gp���X��X���S9=�#���^��*4��ԃ&���1��j���	��>8lY���=�� B(G�?��@!&��C�2`Œ���tXZ@)Ȃ�˸�s���Z%5_T��#Z�jG�G$FTi�r�8��Y_�O(䳅1��{��j�"U�ખ,k8�V��D��P(D��S��yQ��_
6�VVT��w �3Ƴ�$�.�Խ�q��ب��.�7[��g6��S�uV�!<d�oF�Y�������� m	�W#�X4z��o��/8���=]0�/ꘛ?���w\�ֶ֏�>=��Q}��m~f��Ǉ�5�l�o���G���9MD���/�'�fcA����%�����r<p�n	jR��	[���C���	=������k�M[���\�Y,ɸ�(�urB�"��.���?�#z��D��j8/e�%20c���:|`�_��b��'x-O��,��{�d�|nh�5���7e���������]���X�c��AA�xs�%%-]Qlaf��9~P��l)1R��l�媓���VX�4���M���z �O۷2'-X�r�������l/I2o ri=����q�?=�w=n�P����&m�����-��׿*� |���K�@0�ᷙ`��;���;@�9+�U���(L�����G�'1Lj>O�i��n&�%;�~���z �"����,9�Z������󶧽ψ4ҙq��|b9��oN�I�!	$&-��Y��g�U^.h�՟��<u���XlxVHYEB    3927     fc0۶=h P*̋�]n��M����1��L����D��==Z���2�#��	k��x����]�k�� E�=ʖN��a��*؄>ռ�\9bܴ*��Mo~&��3��(���1�ğ�n��ᣃ�M�rS��;a���V"�aYvD��s��l���,��+˴�:��u�~5�1�u�B�vL$�;qT�V���"lj�AXԱ�L���<��uw.���<3��)(WU����<u9*Swr�:�I�e47$�
��Y���.�³���:�p/:����X+�>/Q���\/=')��V�d�$�Q��%^uaC�m�)�Տ𡽾����� -~����2Pq��T���9k�����3&XCg91ѱ�b�`��.N+�
�F�$F��NNv�ɒY=x稦r�=��c�<l���Ὀ�����GpD��Qz�)�<%Y���&è �t���1�!w��ȋ��󗯲w����Z�c���Az������`�i�jC���8�ׂa���_΄��O�[���T������h&���Ô��ŰC�J���<�T�c�r�S��f�=B2 G�����g����t����A��U�I�����?qw�)!$2�z��(u�T��t�J�SA/���D7��r��Rh�ї���l@�j/�9��(��MI�ݩ_�&�RZ�vX�1����$���8���ZY�/ek������G�%���$��ɼ�`T�*�����?}h�;�4�=%g(<<z�2�R�%���O��A(OC�YN�����{�)3W�$n��@���nK2��{Y:|e���.�H��c5H��L�s���BR��B��-��"�}�^�@{B8�5xn����c�Cfw`FZc�� ���$I}!⥅��G�/��N�ro>��u��� c�E�-i�c��|���ESW^��~nȜ��a���#�颌���wq,j^Bn��5�fK�j8{���,C��_����~�����뎢�&~�^�77챀�6c�]��$F�{Qa`;�� �f&#8e�cA���*�s���B�Y6��Q�����v�V&EE���#��l�2�SI�������bG��k�>��;_m����S�=OyS�]�^�[����q¼�B�PC��msM�>Q���Fj	��t`t�D�/_^/!��4���M�sJb�!2���_N��D��i���V�
Ӯr%g.���74������m�� ����
wQ��E��&�mQ�
5$��4�@�	d(`֛�_$t3u$/R�팫+
�)�V��c��p���ꄁ�����]���OT���k3�P,Kq''}�|�UԈ	��ɴe�E�c��;���f4��.�/a�8JZ�x�,�D��i���8�r��m����F��abGo��m;�:����ᖊԇ3�s��{2��x�	�E<D Rh��k����������m=7k�;n���,��p�944�t싹����+ .�E���ph���˃�t@Ԓ�`n̓�Y0��=�Y�3��ܒ��� R��y���{v�� п�V
q�!�+0ҧþ�|4#ߜ.�=��U7���U�>5;��U�|����1��E�� W1H�? !	��X5)�!����3En��v2��hfw����Q�"�m�'5[aZ=��<�Fs�:�ܦI�\/��[�=
ģ�<7�x^�fp�
!��e��k�ˇ��,�3y��Up�Q������Dѝl66Ψv�a�N3̦]]���dQ�ٺ=�h8�r�6��ݾ�%���,��%QzO����e.=�r�p$��,�m] 8�a�Ά��g�d��Bhj���L1������(����}����.��Z��N���)�·�g�:�?q
�H��7]l}�p����#�2
v)=^[u2�/�Ek=F%Ú��z�Y��7�15�)��&:��T%��dc�U6��K18���`�ڋ� �wp�h�Q����V\.>��}��3�lN�3�'�X�������t��y�H�"���-P񵔣�S1����*�]�Ĉo�����f{��%�-Lը@��(�y��EB˴*���͘�ҬL1[�a�����z�m#�I�K�+}��(��z�e:�٨�΋����(�)�]������<��]ʳh��]Ƹ�
��e�K��a^ZA�zྸ��>(&�:E�3Zĩd[u&��J"�-$�'oN��?K������.:ϟ-�F���&0:���r�B�@uł��L������)=�0�,7K��١�N*�{����\�zF��RZ��K���;�PJ+c���P$���h�r��T����]a"r�=�y�=,.����)0�Ȅ_���|�O���JmQ#���y���@[�U]�5lv�K%�H�=�Kˤt��=��/�<ڟp���k�����$V��ܶ�s��F1Od�y�TSh��O}��Y_��ͦݙϤ�= L���]ф8�d1���*����ˌD?I�Љ�Ҩ���P��/�E {L�Fq1�;�[uFoG{�QqtN��p�$%�I�q:�f�\��t���� �� �PgA���J��?�"�K_P��1#E�bY��3�ـj���Q���l���֤�t����P��s)�aZ��ͳu�r�����
9��D_5"\������Λ�>v܇�9�Ļ�行G�����&�otC=�ӊ��}�W�@ig������:�N�fe�Z�w%�<������ڹ���)(h/��K� �IMU�'��ג��?Fo���{kER�po��~�mW��.[�z^;�	&��ކkl�`�T+��9�j'��ց�����Fy� >����,�N?T�i�m;̸ �!���z#���H���O���e�M����䗭�L�MB��<�'BN��sݖ��{����4硴߻����[�,��C�nU@��.�F�\RsY�#�O�ސ�YG����e�E��є ���B�p����6��vniPF����|�E�HA�������TP�
x��37�v�,/9�%9ͫ�ՆB��㑷�A�����Q`2>���.z,	����}����^f�"�fN�{��Ar�*��,%�ҡ�^O%,#X�p��O�>����鞏K�`��L�������`�$�8A� ����*B���X��@9�(����mPL���"9�9e�+q��[���h{���cx���N��k͈���|� ���g�:�v	q�����ݭ�tXVQ)�m�{���j�}&��,	<��k��4=)Dݱ�����A���9���|1E��b`��֦\�U�<���>���L��KɊL��`��XN_���Cx8o�)��ZN£1E�#�k{�W�����gY�W��(S��z��ߌ�7BZ<f]� �ǣ���� Oiq��屫@���h'ItӲ-�y�m�^��lI{��������R�X��z�B#��W�կх�z�͗�]YW��˛�V�1b�.�ʀ�u紞n&p!�g��XFI�0�{c�2�e+���e!n�G-�� :�h���k��5�R�N�uy��s>��%�Ҝ�d�3f���w8ڌ�}���)GQ��t�L]���K<=�4��Q����]���Xqɰe;]ژ�km�����������Nc.d��"�;��ȣ�[=��A�h�LVfdG
#��ڛ�+*CQbU�mF%ĎD�� ����w��W��!�];�nmv��BQ�n��۽�C��rz6W��v_2D�2f*���������3�@�@��P�\�^/j�௓�4�������iT5bJ81R������%@3L�|6F싁���.���
U�%/y�B=���A�G�Hh<nS��Xd��M|���NL��u��+D��� N,�z��9t%��wO5B��H2�`�[��>�MzB���� �0�Qؕ����2#M�tW�X��ݔ�+: �1OPZ\,�x(�����ӓ?�z��ᨅ�7I������ߛ�