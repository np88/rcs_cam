XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��$�!(KN�]�P%Ia�gF�3�:�/CEB� ͅ��Mt�c���s�����]�|�ipx5�����Ú�W�q �k�+j�#p�ș8��A���ѫ����ݏ�D��Z�8ɗ���HbqL���'���|d�{����!�ol;5�8FҪ(�gG�P�E�r���'ބyۅ�����j�Ŕ��׼���gQv0$Grl�%�0�}jy�����ᢢ���,j�E��$Z��ԍ<e��L��B�<�\�nU�X�م\��Jj^FL��O�����#h<�B& 6�Z�$='6d�hH��,�"�]:���n9c�৭ !6�4�����5�>V��W�
v�_�Q:dW�G���N���?�������ק��q\H��Z	� Ғ��m�ׄv��ڎ�ժ�!y�
����A�{pU[VW�ڏMZ��ʢq' ����o�e����ms��/�'�8�q�\�Dyҵ=G�Jg9����ي}�
�4O+���j�(�ҳ�2_�K��� �{J���w\�y��C>�Wy�+hG�]���ƿ�o�G�̅1{Y#���}��6H~����������䱳#m�u�悒����*��
��t9��&�_]�����DV��R�V��\�^gGP�2��\����D:��2q��/1�Wx0X'�Qq�V��y�q; i۳[��|^U#b�̝mZ^���v�5Z��y��F���=����'�`��'DA�X,'5.݊�/:���UXlxVHYEB    17c1     810!�sB'��%�v_���?�1qi�%XW��w_��0�����h/YeI�ċ�d~��B��Ŕ�dXS��`�g=uOM����jFL���Eư[��<ޘ~�%&�'J�vn|��-���?���������G���\� +�ٶ)x�^\��2�ؾ5,����e���=����s8��<Ukg���[�nD��c���1���sv�ޢ��s<3��"|El�:�3�ky0\�ϡ]��[Q󶜵.�0�z��j��|c��[���R7�g�)�����6hG{8q��d����+SL����^���Y!���(s����d��7I�x4���4��mH)
Heu��}\"�n2��]l\��}lSI�����7�Z�{�Ib�P��=��#��$��I=H>�ɼ`�i��Q�n��Y9����5����*P_���c�	%��a_KZ5���x��?���߮աabR�5��/Wx��#b��q�:�-����bwΖq.�6���ڢ2S����"Ą�	~uKi�M���o��J�Qn0����N��l��@�cs�&�])�T�b��ܘ'+�6(�3 YE?=%:�M��<õ��J��Ѯ�y )-���L�H`.���qh��	��������f4��*��+�G�'=���U{Ѷ- �F�s��f��Dw��K@*�l��'�G�y�S��!�^}�*B���]`�dY�H��|�Vξ=�������u���p��el�잙�Uwx�i�/H�?1��G9SW�v�������=�뢔Ng �k-A��E_M��%��${h���dMG��Ү������)��?j�eBNk��g����W	ˈsUvh�\B�)^�YFEJ:s�&4�;���,�$i�*�i�#Ԟ�4��;V	�������C��*+�f��C�xjg�_\��9/!A~���_��y�P�]MPC���U`c%�b��҅�v�us����3�J@AJ��=L��Q�$�n��"#p���ʌi���^n�4��a� 
��GC�"�}b���.�Kʍ����^�3��S�h�1�,�-,i�R-b���ج41�/�����N���9NZ{BN��xVws��8�8Yn��S*v���	�ъ�k)���.��_�}��7+>��4bI����9�@��g��P����y�B7��'S/�1T�]c�B��KƼ�H��씰8'�Iz�4��o�5����So�����2�0��%ɷP���R���P�0�٨ِ�ާ%�;�>��%�?U5v%�� 2k�:l�L4m*�GFp�4�u Xg�'$�sC�Ŗ*��~E�N���8��zv�K�+q�@���k�>N�z��3v��I򋞭mg�Z&����>�����S�%�'����v���)�����}9���Z�P���WM����bi�1M�/15�W���j�,�^G2#���[�f�~��(w���+~r>"mABzt�7���Ⱥ�%d�j�V�jݙ��E��NbG'kO������b�jW㒃NKv�ܒo-��KN�A�R��x#FCE0�,=y]�@Sq:3�XE��_ʧ����UY��|r���ɣ��P�x��v��<'�j�a %�����,ݣ`��0�\������M:#�l ����Kl���l҂_�B2Q�ÄB��$�J']����B�x�X��E���{/�Jq4�S�^l���Ao�-��y������֞���Yf�)0��"Bz!���:��Ѳ�sW���_z�ͥ��1
����s��U���"n:c�K�g1�/NujY��l��?�$}s��+|�a|
Br�h��oF<o��.��s$�|H^�2�Dm���g�A|/��ҎΉW�����d�Uֽ�{����";���[+IlDUA|�~^�t^7�H���8�����Ou�����Npπ���%U�6!R��V�~���N������{�YI�(�X������:�S�j'1OSfc-�GH�A�DP�T6?�F��7����J/C^�L�w� �Ik�N��EfeFxPN21Գ��s����n�?�df�