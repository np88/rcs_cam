LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MB IS
PORT (
	fpga_0_DDR2_SDRAM_DDR2_Clk_pin : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
	fpga_0_DDR2_SDRAM_DDR2_Clk_n_pin : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
	fpga_0_DDR2_SDRAM_DDR2_CE_pin : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
	fpga_0_DDR2_SDRAM_DDR2_CS_n_pin : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
	fpga_0_DDR2_SDRAM_DDR2_ODT_pin : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
	fpga_0_DDR2_SDRAM_DDR2_RAS_n_pin : OUT STD_LOGIC;
	fpga_0_DDR2_SDRAM_DDR2_CAS_n_pin : OUT STD_LOGIC;
	fpga_0_DDR2_SDRAM_DDR2_WE_n_pin : OUT STD_LOGIC;
	fpga_0_DDR2_SDRAM_DDR2_BankAddr_pin : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
	fpga_0_DDR2_SDRAM_DDR2_Addr_pin : OUT STD_LOGIC_VECTOR(12 DOWNTO 0);
	fpga_0_DDR2_SDRAM_DDR2_DQ_pin : INOUT STD_LOGIC_VECTOR(63 DOWNTO 0);
	fpga_0_DDR2_SDRAM_DDR2_DM_pin : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	fpga_0_DDR2_SDRAM_DDR2_DQS_pin : INOUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	fpga_0_DDR2_SDRAM_DDR2_DQS_n_pin : INOUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	fpga_0_clk_1_sys_clk_pin : IN STD_LOGIC;
	fpga_0_rst_1_sys_rst_pin : IN STD_LOGIC;
	gpio_FIFO_almost_full_I : IN STD_LOGIC;
	Push_Buttons_5Bit_GPIO_IO_I_pin : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
	gpio_FIFO_rd_wr_en_O : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
	xps_FIFO_cam_data_I : IN STD_LOGIC;
	xps_FIFO_data_rd_cnt_I : IN STD_LOGIC_VECTOR(0 TO 19);
	read_clk_fifo_O : OUT STD_LOGIC;
	xps_epc_0_PRH_Data_I_pin : IN STD_LOGIC_VECTOR(0 TO 31);
	xps_epc_0_PRH_CS_n_pin : OUT STD_LOGIC;
	xps_epc_0_PRH_Rdy_pin : IN STD_LOGIC;
	xps_epc_0_PRH_Rst_pin : IN STD_LOGIC;
	DDR2_SDRAM_VFBC2_Cmd_Clk_pin : IN STD_LOGIC;
	DDR2_SDRAM_VFBC2_Cmd_Reset_pin : IN STD_LOGIC;
	DDR2_SDRAM_VFBC2_Cmd_Data_pin : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	DDR2_SDRAM_VFBC2_Cmd_Write_pin : IN STD_LOGIC;
	DDR2_SDRAM_VFBC2_Cmd_End_pin : IN STD_LOGIC;
	DDR2_SDRAM_VFBC2_Cmd_Full_pin : OUT STD_LOGIC;
	DDR2_SDRAM_VFBC2_Cmd_Almost_Full_pin : OUT STD_LOGIC;
	DDR2_SDRAM_VFBC2_Cmd_Idle_pin : OUT STD_LOGIC;
	DDR2_SDRAM_VFBC2_Wd_Clk_pin : IN STD_LOGIC;
	DDR2_SDRAM_VFBC2_Wd_Reset_pin : IN STD_LOGIC;
	DDR2_SDRAM_VFBC2_Wd_Write_pin : IN STD_LOGIC;
	DDR2_SDRAM_VFBC2_Wd_End_Burst_pin : IN STD_LOGIC;
	DDR2_SDRAM_VFBC2_Wd_Flush_pin : IN STD_LOGIC;
	DDR2_SDRAM_VFBC2_Wd_Data_pin : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	DDR2_SDRAM_VFBC2_Wd_Data_BE_pin : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	DDR2_SDRAM_VFBC2_Wd_Full_pin : OUT STD_LOGIC;
	DDR2_SDRAM_VFBC2_Wd_Almost_Full_pin : OUT STD_LOGIC;
	DDR2_SDRAM_VFBC2_Rd_Clk_pin : IN STD_LOGIC;
	DDR2_SDRAM_VFBC2_Rd_Reset_pin : IN STD_LOGIC;
	DDR2_SDRAM_VFBC2_Rd_Read_pin : IN STD_LOGIC;
	DDR2_SDRAM_VFBC2_Rd_End_Burst_pin : IN STD_LOGIC;
	DDR2_SDRAM_VFBC2_Rd_Flush_pin : IN STD_LOGIC;
	DDR2_SDRAM_VFBC2_Rd_Data_pin : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
	DDR2_SDRAM_VFBC2_Rd_Empty_pin : OUT STD_LOGIC;
	DDR2_SDRAM_VFBC2_Rd_Almost_Empty_pin : OUT STD_LOGIC
	);
END MB;

ARCHITECTURE STRUCTURE OF MB IS

BEGIN
END ARCHITECTURE STRUCTURE;
