XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��i��~����aV��Ox��*������@S�
q���)ГnZ�p(��''���^o�d���M�<eޥ�F �d�<�TG��(K�>q�+�q(LL%Kw���@��T>ݬJ�������R-�t�s�T��,�x��2�03f1v�l�ŝ(2�x���y'��`�u�1��^8@��E�V�h�hC�yM]�r0UYG+I����e:��N�,�t�7���>H���*�^���,As2?VV�7G?�e��P�]`"ĉ��ݮd!�f�����*��?n�tă33,��Q�5�I���:ҌȺ����o׻�E�)����Z���#+�s�֊Y^�$	�L�V��ZN��b��3�)s���H��{�f�5u*gN�h���#1��/�6�R��]�tt�%�bx�ҫ����%ߑܪR�Q� � �ȊO��!2SK�h�'����M�&U^ħp�	�>��"B���Y��$b��.�۪�_6���gG=��$���x�A��,P��|��9�FQ���6��l��L�m4n�r��f�H�E$6ӻ\�E�Ӡ�\�8�N�=�_���.���`*:�|3�!����-ٰ<��ɦ��5F�A>٧�-�U;)x�꼰�y=�d�.l�w�v�b���Z��ӝ�����:6��聓b�H�]�����N�r�Æ�0k̕<�^m41� ф�:�1_w���Xv_��C�q��|:䝟���9C��;�HW��GJ�]"�W�=�os&�+-x9� FXlxVHYEB    507a     f30��9��qkǘfF���n����j��gzss�E8������D`�6ި7n� N;\�可�IV;B�:�jzVx��J��,a(�f��vv�$n�+�c._\k.۲��u�����P�js#X�eN���X�QqS��R�����1o�ޮ��&�ָ��fo��#6]�o�V�S {{�l.���~f�˖$ �(�"j@!4�h���d�R{��9��6�,�������V*Cp�}ˤsR�r�\�9��-��¦���W�z�	�a|�
O2����x�0�h�,(�7�g5� ��'�����c�Aʣ4�e��b�=��c���x��{ٛ92-���e��������5���(�v��Ky�eܟ7�=�Eb_ǒZ���
1���лK����3kV<Q�1�.�ਦ��c�v&�A��f0��if]��^�$�����*F/�s�&y��|���|�T�v���85q哨=+�L��������Y�A��>D���+��vV�pw���$�-�P���6�Y�����f��c{��[ֿ��0~=�Ҋ���2�o}���$
A�Cȹ�.�� ۊ��Z+���T[q����O{|z��hP����JV���qT�<�X��T3N�X
��,�LS��sU�j�q]�'�}��p����@�/���)�W��E-�o5��-V�)��������L�YؼY	�ȅe�����(?A}U�x�XS�w4]�����P��%�ne�&� �^2)��pԛ8���
l�P($rQ�����j��~�0������|k{;槗�W��P?���b���3��K�{��E=�ƫb��&t�	�3���#\�w���y2ᗰ�}fO~3����D���>���ޣB*�[��u>M��E��)8^��� �����|�U��,�Us�;N�#�MYI����6��~3d�5R� ��5��,��[N8��[Bx����p��s`1k a�I�]�x�0�Qk�bfI��%�E�E&:0a��:�ڧ,���������?/�t�[|��:�Hx�$f�'���	'�)�bC�#d�}�Kkӄ-�@�y"�v���%�d~��N���r���ᾞ��~�����h�2ꇵ�����˹ڼy9��F�
�6�3z
��K�n��45��V�[=]]�w�"cI"vSB��:��ͧ���S8;'�9p�0��dJuxI��P %3��{�;��M�ڗ-$���,:����*'	t�� �����E7�	+3��u8���/�m4
�"��;)FI4�>e%�AG�P��:G�?G��ČLv�þ_�N&���~U@��W:�g�._�4e��T����[������
7%��i���C��ӂr��ek�˸��"ײ�Sr�/í��
琋�H��S�&��/M��$�Ļ{7iɠ
S�R�vh���Z�Aז�=A�@,� s2hE�~��:d[�1���'��rb��#3I't��]�_39/繭��,T��p�������4�vs9e��ܘ�^Sd����nV�e�T�{*�-^t7'���ʃ�^|"��ywI��۶� �;o�h�E�jö|�W0����=5�ڝazђR|eɦ{z�=�Nܜ�*r�2$A/�4ST�.��eb�G�����%15������?��Lw�B�%^x�E��?����(7K<\�b(ܥ��ۆn���+z8>�lE_��!j��*�69Ѫ���wW�'����
����^Z��Լ��7�kP��)����k("��}�{u)�z(�58Q�Cx���6�5|�+�~�tn'7W5��>�][״a���z����Z������8L�����p]Iv�.B�D�,\:J�.kQ"��["�Z��ب2�ެ\�H��O����]��v}T����0T4�T��N"�gAt�ˤͦk����`����}?���ee��AZ|P��YM�b�a�T��\�]�t(.���c�}�T����ߴ�r�4*y� %�{��x��OZtn�h����1,��ZXT��K�u��������#"��Cjǋ���*�����z5���S��*��+��.� ��"�;`�lǇ���n-�/п<���곚u�g%��ߺ-�L+�4/`Ѻv�g�t}w���}�6Y���W�ތ>���2��;K���(���{MV�oO��X��'�xZ����5+�����P{�r�H�5�=#X:L-*Ђ$�!�@��,�VИ� �2�|1iO�o �o�8ن�:j�r�3�y���V,�c�&Rn��d�4�I>���&��?�l�j���B��A\T�hA���K&�� ��=M?X>���=���ȿy��L�5q������B{6ɽ"'7�'B�
��b1.*�s����bRs����<䀿�Ծ��F�{3~���?&�a��l�	�>8#�8wn3�����?vdjH����ƃs�&��WҰ��8-���x��/c�	@ l�l-8S�P]~d�����?��!�l�Ȩ���;����A�۾�b�kS@
�"Rg~���3�u+�g��|zٕ� &^%���x��'!�%: H��۶p�ݜ걿[@�]<�%o.$u�mK9��^���v|>�k�T`p�?�X�"PM2���������ɍ��k✸֔c)���"~�C���^�@�Ȼ]������	�B���g�ى"���
���Ky ��w/�$��\�u��_�~{�{5ثb�5��I⡟��~��o"�i^��4�=.X����*�-ͨ�Z�Pٔ�M���}S�G�j��Rd.�'5�N	��������O�{��dX�]�Y�MX�]� �_����L؀_n�o�O����)��:���
�HX���{� �ʸ�����J��Q���vxT�*���dr9'���b�vj<`<lFN]�S3B��̃��M���'B��� ^d�H�������]�a����pf�e���`��3�Z�A��TC�X��I��:�|AȊ@�,���[�g���c |ts�?��]�%<�d�NP��(��:��4��ٵ��z ��<�\<��� ��O�L�<��dтmZ�G苜w��Ǝ�އ8�x��TY-�2�i;�)7�V�|��p�\�$.Sq�m�����Y�	��ryZ)k�1��c�o2�eA����g�ž�[K�僎�a>�؀��/�T�4�i�V\V~�@��0[X2��1���:=Q��w}��|pc�VB�n����s����2Z���z���k���
�g.����G�����d��-��kf	7`�N�ﳝ[����%Hi-Ȁr&JW�Z�MG��0�W���g��v�������l:�Fu���ȗ+B~�Tf�v�e��9sn8��鬷I{�#SM�8��5�*����7U?�܊B6�b��Yx�l>��_�f�̍n�r.%w�6��1�5��:ְ�|�n�o;,��PϦ�I�i2�������{���|@gCG��^���t�)Mzϑ�e���P��sk���Zt�aE$��q�B�J: h๶��z	�kS�臘���Ά(���C�G���=_Q-%�Tc(��!�=2�-G�\����/ؘ�λ�W�Ө�U{PP$V�*R g�9(��N��m]���d8|Qz���\�x�v���ß��l��g蔒��[(]���B�Ǿ���^���9�����ڟ7��Sx���T�h�������كZ��{�;���s��r��w��[N�l ��+	��X���_�܄N�Ԫ ��S�N%	h��9�ع�Sh��,)[�BYq�%8)�+�p��=��s"hb��q#��]�u���͓a��9�^�����/�:��g����/�n�JQ@ҥ��.���