XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��M�;�o��U$r������ߪ7�k�gw�۔im2VY�u�т:�!nE�(zdW��Cʍ��m��V<�������{�H�������	��7ޛ��-��H�~������/:�hƠBޥ(�q��T����P�u^�zl���@�J�[r�NI��_Yw��8�v"�����J��w7�%��c�@-��*�8.4w�J"�a�l ������7����U��KB�%a^�.���h
�HKZ5G��4�7���`AONv���=�K��v�ɔ���v����dP%֣��fh0.�i�@.�]"+�V=/n�߇�/7`v������O���{a����`9���T����DW��� o�[UY�����t���ҒTR��d����F��=�!A.�
;�Ç"����t��ī�������Rh,�%��a�'�s!���;Ӧ�<��@ؾ���.��4]�[����(*1Dߚ^9�����E�}f�5.֯�1��6�m�w�c=�S^�ۉT��m�Ҥ��t�tO�����@���H�[%�Nk����(���[sōkո6��[a���o6�Sk[F�5�aKĳ+yI:FE �y�e� r%o���2���q�K$��/���]�:�餎�9��k�LT��&����{�/�EC�"-��$jc"���b��Ԅf���K�	�u2e{��k��Y�pC�0���eꏠj{Fk����� '�O� ��؞���
i��m<Z#ܜ��8�\ci���p}d~�x�2�XlxVHYEB    1da6     940j}��I�	~�FQnK�tC۴y]��qc���ǁe��h�[�a�
@n�wS`nn��~X%��Oxi�f!B���F�A�]\�/�B�霋�#(M���������хҸ/&��nNK��i/�4�܇�U�6�ەf#��NJ��*7G�Ǽ,������^�8a����&��a��S�{N=:�o#!XxR�LKS�B���9����-����y��4�fHU�h�W�,�H\츠{��ȱ�T�`��H��8n*�oD���gS������L�|���9_���L�V�!�<��-M\1^츉k:�UJև�~��w�EHD�4u(~���%!uq�4x��EV��bXea�]"˷w#cܖ��j�#�gߕ�/¡��q�y:i-xe�x#�9��=ϲ��G���ƌ�u,и�i,�ܚ���G��K�Q���h���T >��>�	Z-�E-�E,�)[g��$�V<w��b
j�&�	*�88Adg���d�Ql��7��M�N�����v��.�yWU̝��}����+C�HӋX\�J���s5��yR��gT!QU��S4x�2�oX:�K�Z�a?�;�WU��>�ԩi�m�]�m��Rd�q>\��_׎|���~�Ζ��'��\[����<��="��s� R��B����w��n�b햸�x�l������=��ݿ��msB>�*zc���鞥G�3z
�\ڮkP��L�*k�͋��&���`ŕ�� ��U2s$�.ݱ`�Őy��@Ϊ�x?�f]puk�H�R	_jg���"g�d?1��%�3z��a���s����Q-9^%�ٞ�� ��D7H^	��QʃmՂ��8˦�>��l�&�p"z�}� �>J]4Ro5���8F�1�a�@�vOȱ����=����\d������&����*�2RL�t��B���,v�=b�'���n3I6�T�p�����\~<�����0S� �đr�6���x�����`��S����2��ֈI�'p�r��̵�oc����$V�]s�a�t9�c.�"wsIЍ�����#�
z޻̄�E�P�8�p1!3o����9rzE�-��m��٫>'���Ό-��q���K9�l}9��Ԅ��1�>�B/�1ZǏ����X��$��k�ݛ�G�ll�;��eF�ߋ��^W���F���)�X@�`('
�`���t���x����� 1�)M��i�� =�`Ö�i��RI;�Ɠ�u���Y�jڥ��`�e��Q�%�A%M1�Ċ�5�棠 �9��!�霸�?���5�^�{�ke�tuO���H����"B��Gb+�"YE`}�Dj*���(�����Q|PP�1.V��h���V�l8�`��I�B��G�w;ʮVzܴ�;�UDT/�!T���B��k~�Y����Z�ͰȆ0q)��i�F0
�q���$�K�o��f�ac�e�Vmtm�k ��1���/�Z�6����{/�]�WД��������j�A*P�0���5G�^̀D|g�gjq���j���(\2���H
_`	8V��{�/�#��ݐ����G�_u�T�tgq��7��V�=�fmVq%h���5�b�;ڱ5�Ȫ-�i@c��	�/Ơyo����Yd�m[*���~��}���2+$�_L�~S6&�Ͷ�������@.	煄_X�������t�P��x�B�U[��*��=��BF	�Q�H�2���0�(n[`^'��j��Dd���򱡊�}�,�C��pc�'͛����?����6 �sa��u0��ǎ� �u�J�3� ����lA��,>�=�G�����G��~��'���m������ɡ�Zk�I��UQ5h�9�"�L��6Xй��2t���9�zk�E4Ķ���Br-=��[qi�ʅڌQ� �m˦�l����@�9��<�TF`���؇W��ʔ�vK��5$)ò}{��P;,8�@�P���#���9��bf�ZjxO�>|C�
���`65���,
~��>\�Y!o4����Qf�":Ը/l�)��<f�]��ߏ������/����φ<3t���imr����$�߮0���b$^}� @b�Jr��y�2�U#��e� ق�U����*E��q��<�>�'C�/-��X(�q�c\��j,�	-�Z�:�P/�
�{�>/h3	��ʍ�U��~�NITHZ&{GDi���U~��Z�6�.O���є�A��o�K�A�yI֊Ч_3���i�BDB�nU�F��p��������g�W� gC(&����n9��c�b`��/����"q�E����Q�����v����JJ��K�.��g1�3VE�	:���dp