XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��gM���Ӗm���ЎE-� u��y��3�6AY&wfSQ����%�,'9Uo�u�� ���}:�_��7o����0�E%����)�Ne�֊I�x��v'�FX�p-��н�D2�G�=.�>A߹T�;���~��=��}��A��]��D[�œ�be6m4��q�{��q�3�1��۟��;�	�jRɩNw���fAC5�܎ ���C�mM��˧�ݫ�)\�"�'w�),;�X6&�\���1r���kut�����b��	�}�}&/�]τ By�����F���m�����E�>SX)+���Cq-���	,�G�mW��x������<v��y�S�������_�Bn �P��9y�P�[N<��R�l�XX^X�c���t�Ba6;䙏�X~��	�l�%g����&]�Q]�<]}5+�/���QI(s>�Iu��65�϶g�:d��Z�cw�p1,��R�9@�
��O�����X�l�FE�D�&=���{-��Z�|��e?�m��l�֣�(�fWI"O�%ɻ;.��˧yT	@�*��x��KC��%Zr�� 	���.L@R,xayk`+�A�����)��Fy��r_�F�wJ_���`-�2�f�V���|�G���O�J_�,c4sD��>��"��Vu��XK�Àn��Gq�a�H�]�.V4�;|<
�� ��D���N ���:�F4�d�m�؄Ѓ�0J����L�]�6��X�Y�^	XlxVHYEB    fa00    1fd0�w��wG�I�ZS�E�F"Q2�۟�$�n+��z ��ط}:s��{��=��Wf��e5Q^ˤAx�,Қ�*E� �m{w&��Y�l�&�V����U�,�Zy���̋R�-]2��W�?t��2�>���]�{�1���2�����5�95�92����<ɪd�������B*ڍ�歶_�19��<Uq��aEŏ��ݑv�)�*��Q�+�Rx�8+�b*�(��+���7ZV�O��#0�5�~��*�M���?I8�k
od��s�Pj7[�� $b���<��G�L}��׹ؘ�W?d�Ŵ4�L+c��A�R�7@X�$>��3�'RF;����3yx��#X�Go���v��{�����ګNF4q:F��iX.\�o�n���*Td���U_��	pgS6��@^�Qk��b��)�2�p��j q ��e���{j8��t�?u7�U��ottm�B������.�1ro���E��DT@���4�"���אX�V;��4��k�zu���[S��7qO�P����Z$)�  ��I�	f7��yQ綒�/٭.�'JX#�>l�[<"]B1����fg���B�l.���="2�6��&V�d^d��J��Tti	��-c��E� �;e�'��%��aG�u�N�/�'B��Ɔ��$dV�,�%��&���9M�Jm��4.�|�D��i�/�e)�w���oqÅ �J���̰S�1�t,v�N!p)n�G�������_/���/�Z���>SB��+����5�:+(�����C̬2^'_m^c�5�?�U3�����P�LR
�?��ua��Մ��/�,�$��5[�(����c�KW��O�V���*��T ���쎸yy}Nf���$y����$Ʃ_��Ot��N������<����ޛ]�E�޵��W+U�f�H�2���V;[A?'iI,����eN��.��E��Y��������c�ϔ�+� ��
�ꜣ/�oՉ��"�º�jʹ��-R�T �2�6�B�$�n�b������{�ԏ�!0(:���-�jږm�͕�Z���V�P~w>tw�mbU��W/�l7>5�fz2^��X��~V���䄓t6O�9vx|�����	�A����$R�!$F�*\
�2�ek6�
���Ց�7�xO�b�~x��qܡFj��B��+fNE\��!���>���X��f}�8V�xا\��/�l$�F��Ȃ�G4��=�Y��R����{�HT��"#���������~F���������sٍfڔ?��~�.�Z��(���(6���k%rS�.ް�"�0H]�]�cy˵~Y�WkY>{�	夶n>@��q+]W���Oܖ����X
N:�c�S���kɭ�����w5�o�~���(z�j["s㹫bP��f�۫���!ȍ̈��e ?�;y[���kmؙV���i�~; �R�#-�r캃�,�RH>�V5�"_q~�tJC<w�i���a�'ۮ��kmF��p��&SwR���P��������FϾ� 3�7B]����"�6�7�F�l��84�g�Q~1�2�H���MѶ��A:f𞃹�*�e��c)�#%J�X?�zq��-,����0k����S�"���GR���>�r��g6E�.L7x��Q�2-|���mf����V$=��0�Vd/���6��>C�%�Xp�ǁ_YǹQҖ����?�+ަh�r�;��Ĵ��wHFTg�-$�F��F�-[�rbZf����d1$��2�X�}��-��|'�zu��xó��=���;~8��02���r@r��l�ż���Z�I2GDA�H���ٺ������Z2��lU�a�pF���!���h�;��61�;�ly)��Z��Zcx�g,+���jM$�,��ǏI�F7^m�bs½���No�>����zzrV\	p��ï��}U�!ǳ� �?��Y��󭨖�h�9��N���������[u!dޏ%c`J��T�}��d,s��n@�˟���Z�*��P`���cR��p[y�cr��Z��FJȿ�4��F�y�U�P��A����M��9O~�ɉe_*�XON�@����Q�i�,� �L �t��r^޵[��+P�'�!���v>^&�O���������&���\�,��_�Q��+a����ٰ3U{(��"�')<z8��e��Z�jh	��_ N����׶��%⍿%���T�#�{���6��ȩ�c8�E���`�V���f\�(~?�]���d�GU�<���8<�b�O��/���
w�Y���Ұ����R��Zn\<��*�
��Bw���4`Jy��^L+�iNs�dr7=͙�����1Y��)����m��#�I���0s���'A�H#�GM+GX�L��|��y	[}�W�Z`�J��_C`�dJ��3�v�&���`��;s%|��3B�Sh�A�a��G�n zy-�D[e$�Y����AO�5S���,�3������gl?ͽ����{%�Z@����?�{�}nbڶ�A\�zyT��6C&E �f�y��k��U`���'�qXZ���(M���{�̀cLFШ�D4�!^$���!���9)��'UC(���#���h<#W�Lɐ/�ڵ���O���9$��D���G�ϦÓ��)yK�ʺ�T�Kϡ5X`~�3�e�"��=E��!�x¬/�O]�K�S���(<�2�\����"xM����Y[��Q �{���L՞"36=�/i���D�5cm��@��AU��0|�=@.��U�����������k�p���)A���ӉH�&��n�]��ad8)�L�KfvԦ�x &��+K�@yd�U)��~��oW�Xum��%�M�Y���T5tѢfL��M�i#��BK��h0���zN�5���>𢭂�+�	غ_o�>��[��#��Q~�W�&7K����>�A�w|�s�6�T��[��ս\F�*�S*:��ы�� BZg��5g�n��6TCZ�����N��9k��]n��P���P#0G��s�_�ת���O���R$�x;���?�e�X�7j�R}a?�qH��K�a�j��]���;����Q�UL/h���Ί�xl�U{��WK3�hH�<f�m������Λ��v5���g1��90썇#�' B�ZC�\Vd��a���ϐ��1	ĎI�꧆���˴�U(�i��u|za��4} �JUq`�ٚ�+ܯm�o��3���
��\���[�LE$����D��#��ω
�ҡU䣷�G���xX>B�sT��3M��	��`l@��1E|��_�qf�~���r橒+g˥תپ�C� >-z���C�	A e-�t�s5$`�f�7[_X-�䂗t�ǁ���T�y=���9"	��e�>32Tk�t�6�j�Q�/��QZ0��O���� h�/	���}�k�;�w$��y��A)�I�N�G��!�h�p�ώ�����P��� ?��6[����M<�� �=�<��OT�ã��U���ү� � z����%U}��!iZ�M��D$"Q�@��g��1�.6N���5j�W3������?m���#�2�.�խ��I��AhzGX��t���?e5L3@����.:��'���Ώx:��#�4�j���kMJ�"��z ��r
�ܯ�=Yc;���`��_Q-&��
��4�Ys{s!/��9g(}\� ��Ѻ��+�D���]�����f#B��+]¹�P��iȿ�C9S��stJeW0d m���,�	��o����������~��_`����M����`T��P����A�=쀶�3
^B3��d�)���Bxfa%�Qh� ���TxY�2^4"�c|��k����G V����'m����"ʚ/�8d���ш�ĥ��+��-���S����:[lS�1z�n�3�dy7�85�o=�MW�j)��C�N�kf%.S1y�2��'�@�/�s�{��r�~�.k� v��vX��A���:�q�O]���(��fUDa`P������<$�9B|��.���S`޴;�S��*�B`�����\,R�� a��r?O���|u��t���+��i/0�~����k�ms�N�������Yo�*�^0�q��6�(u��U��n�}����/?l�R�CÉ�v���K�&���k��F��n��E���j��>P|�{�o�sm%�o��ʻ���c�'"o�#�Y�[rT��^eK*��K�~� U�:נU�ػf�985��� Z*��(��I����ؙ�!5M���W�~�%��{	B���~��W�K��I�8c�;���9�?2����.*�x�u�:�51��Yt�W����I &C�׵Y�P�\��t�}|Td9�����E>�K�|�(�_�GBޅ<�B��	��TC@�Y�@�4�3��1��0m��c') mְ��Q���
���a-�sтt��7��)�g���̈������sm���r��u�w�\L}��/�r~|����g|�����<=~x��O�3^����x�(ll����S��3��r��[!��CK~߱�QBSf��ߖ����	�˳����I_�Z9��p$*O�A,����Rx��$L���AR�,�9C��f�z���΀y����6�b��؃�^{\V6�W$9�@���Y6o|fO�qp���r�ޏ[sf 7���^kr/υ�n�TB+b�+K$�(�Z��e &����	��Y¥�A#T��#�k��ƿ���E@��9/�0�|UEO���e�a��r��d��)tѽd�Mw��#�s�Z�M_���B��W��9��m��B��zx8�=V�"Ӹ�}�����>�#b�($���@��۶ѫ8�X�ZD#c�%��Z�=�Scc� ]��75��Z������r;AYݺU���){Ծ��[ʰ���{B#oW0�^��jl"0fg4��r��$ɲ,n]lA��l�,��#p�es�v��l��9t. [�R��K8/ֽ+#�c0���F��ٛ1�qyв���x҃ݻ8�5V��Ji����Ke>_�_ 2�+<q!�7r�-�\��W�@4�u1K�!)l@e$-Gw�,>��|����rl���O���{�ZG�:�:�"��E�Sj7&$���֢�k���-Z���!Ko�Exd�{��W�����M��_k�
��!X�X;�fz��)� +�hkێ|��u���t�_��Nx�H*0wK�3���'�Ћ�?6:�����q���/��E��ci[t���kp��}f�j�f�n�� ~�H��/�`
9�Dl��>�����4>,k�.�����m�k?��dx1�ER^k.��טH4���o��&��7�=渧���ez��NSݴ9�~B�Qc�Z�l�8�i�����5_���1m�����G�Uػ�"���k��<g'B����*H��P�����XX����@��=�w8���8�����b�LgSC^�r���īF���R�@h]y�}��w67�]�}�������.��u�!֗��}�����=�	��,ym���9���\��ݝ�`��Èa�4�B�a�hP��
#�CB_g�M��,g2 �W��$Yݾ��?���9�.��v���/���Ҁ���h��l�\=�S�6+']g�"6��p��#��u���c>gV�����F�"��on:F�j{��Z�?�ZX[4$����mg��ú��, ���m��$�4�y��Lpoh�}�5���O�b��������Tf`��ĥ�|n���Yf~nb����!������h"IR�_8��AQZ��r�I���љ�/b<(�X��g&�_�aIe��)3|�C����fD�&�h�T_��z��8�<`���?�W7]�SBF�6�{k�>����o9���'M�/��]�>V���f�~f=Ja{�@r=ڷ*6-��D�2� ߚ�q�B	X��iD��G��W�!��F$ ���:}<���K�Ц�
���J�D�_#����K(���E��S>�?�6�Si���Jm*�5�g'mYz���מL��DN7��X������7�3��z�T���_Gp5�������f^��O�Y�9:�U'
��Φ���Xf�&�:	�oZ�&b]Oc���ߌ�Ή��A��i;�QQ�ed��g`��΅���Vtu��_u�˳�yѯ�9�\W�� =6H��]���҇ă���9K>!�F\�_q1#��
�y�l��r��b�Wo���C��P�˶�۰@�9qF��?�w@�2���
p��J��c+�ƧÂ$�v�gvߨ?é��{!�B	�y���Y�ј�����`����V��H�?*��zd9.��\��u��"�v��0���ġ��e۟P7��nE��댽`|?f8�F�п|�y�Y�.�c^{�ƕ���n���������r0M�}G�@��!�jz��Xν2���t���I�������6d�?X�b�fY�5s3���]�0���Y�LS��n�[�\zW㥪o18�ߞ
P���b�ĕ�9=���2Gs<�V���¸/�X�ٶl�N6t]�B�s���LYv�9!�-$9�~5�����`��s$x��N��Xz���Z�jh)kD�wj���b��2�Ȝ}�����eW'���*����c��G��� �EA7�掸�C�Ë��"
��;*���k�!����}W�u�tş �o�Ҽ�QϮ P�z����d6g��y����f����㜎�[��5;��{WzǼ	������0}v-b�+��̊���d=���5�6%`�R��	K�)d-���N���� C�o��u�n#h�Ml�ъ-i���81~u/m�-@��� G�H���[UA�����2�su+o4�;g�? �@�lt�M�`V��f!��s�0�ܲ1���C��#?����x��׷è�/53%M5	GB$��̉ٯ���@pMt 66
�t�Xr9ߍ/Ȩc5�[h\`DԤ�,��A�����u���bxt�d���o����`���Ӧ��^^�8=`E�˺���z�q)�crCk�4��6qӝ������/aɎU����fld�8��.�v<�~���|	� J�R�M�B�`iR�����ݷ���>͠ˆ\�^��CXoH+j?�G���Dxj�z�U�\I"s)x~y���b�)�a�N��h{![r�{R��a���}��lSXTc#�f!�$l?�����d���g�!}p�3�[ǄFg��&h0{�_�K 2�z3m]g��uv3v��KВ��V�\�s�t�8��=E_3elX�,24�����̒U�SN
m'S\4"q�2a�T�|���
{W��@ r�{�ӘU���7��K�������~^���1��,8ߊ�<éy��0U��ܽ�h��f�����lQ� ����z�����N�G���mA�N��*u����x�F��uq�j�K��K>͵���?ۋ��A�dh`vk��6�d��2
�b�^(�/��n����s;t�%%垿:�Y��_�W�(;	::����*��ҐC|o)�*&
�e��0��^]s�{:�Z��eK�^6O�'���FE��U�z�aNov'W[�0�T�G��. ��b�(���
^�J�Z����`�U$��������ⵅ򕪩R�CFC��8�]��i�o*�%�~AP��i*���x�
�W�ٶ�������/�Q�5�Ѽg#�B2~��W�58��'�(��rsH��Zz<DA��mO\>� �N29@rOt�9��'�`^�%�b�c��/+!��B���#F�z��c�P@���XX�HԻ��+���@)s��މ�8�dx�l���糽�~�Q \��]K����U�5��!��M������=�Ӫ��{�,��N�Z��P&L	�qE�����M�OO��4Q��Y��X XN	#��9��ɳ\���g�B�2J]����*����P{������,� �I����@�P�ڦQ����O�_y�2:�
�u��>e�XlxVHYEB    fa00    1340�Y�Z�`��z��8�@|���=:0�v��:l�v����Sr�nD~c�0�b�}5�U6���:�&�H�H/��v����Ҁ� �ʵ��<�*^5j��p�%ف�.ȆmV���ϊ�u��-�C�!����|��T���#fU
.$U\OηD����٘��ш��U��>`̒��f��;���(E����c��3�^�+\���_H 
w<���?�w�Oeo��h!�(S�'� G�ͥ����Y�\�G�_����i�ʒ��,����U�XԼ]�^������	��/N�^�D�3,�����q��;~��=r���>QXc��&��5ȶ_�X'=��ao� E΅VԠ��Y��_B�����Ρ��΁������ۘ����~4(��kb@R�ʀ�t � ��6�vDYW�:z�?+X~���Q��b	������R�ƇJ S.���5.u	����9�ɰ����j�>9fP�f�d��k���ʭ���Z��z:�xiR�,k�S���d"�P��)��%'����I2����ᜎ�4]�P�N0� W��Y)���YЯ�ym,@O���:��
6cL6�o�����Ĩk�G��DX��k���4���(�v�g�뙀�-� )�!���&C��"���}O7m� �� vC9�![N̴��tD��a{��`�Kq�EM5�Qnb:�|%u
g�SǷp��]�w�$�Yw��JLx t6�6�*|�|��v��3�j�<�z�A�P�xѦ�J�l;��h4Sڪ�`�h+�:�N�6ȢPOy(��H��L���G�ڞwI
h�<�q�?��ѺL�Ī�@g��d�����6�\C���7X��k�ifQ��譊�8��i��#Kj���[q�>D�E��Zر'hɫ��Y�ђH2acޝ�#Z���9��V~G�,��É��K��y����썽�W$��3��u �|<J$:'>+B���>J��M�E��d5JR/�M�Ժ���xd�����1�|a�e�82{n���rs55����EYn���.���S�ҞH���LpD��s�ʩ��%�Gk��m�+��%�O8��3���X��O2�*��c�XS:*b��lnݳ�ǜ�����������n�|� ��ũ߼��|Ҙ�����3�*���b�
'4��V������+Dd�(�.������Կ6=:�-�77t�wȌ9�e�����I��<9��sE�Ə?�h�hVFZ���=�PTy��O�Qo�.<x�܍��^U����ܙ�qX����������@�p�9=�s "��b5F�]!-�f�*��۱�$��O������
���s+��D���FT*OT�G�8����֫�A�{��x��Z��4q���V��+��y�[���@�t�I���!�����u/�;l._�MF�Xjn�O��_�lj����@x�����#,�	����cǕ�����C���mh�������;k�.� ��	7�F_�� Y贫��E���J�55[���fig�bl�w5�N7���0e�w#H:�!�6���U5�2Q6����Dlȵ���66�٩>���<t��Pl�X^8M���}�6F|W���gs%�Ȕ-"J�źo2��L��r�SF�U��2�t��`��'<�.��Y�>imY���[6D!�\ �B,X��5�!s���ݠ�B��.N�?���y�ZT#u��w&Ū��{A)?ű}8�2=ib	{�*\k6�H�k����,_l~zA��fv�J
�%-��,N�FZ�1¹�7GB~x"�$�-)Qw���+>�����f�ze�#����,L{F�M�4K�^��5��Y�wt�9������]��v��4I-�q�A�	��}��H�����e�D<�ƽ���@J����a�{����YO#JS��Q�D�橭^va�3&���aW�~&szS�v���Ev������a�̸=���@������2Ôt(j~{V����\c1�}Io<��_�Ք���F��P�a-���$������i���0�Jd��������K��܄<e�����+"�U6�a,/���Y	���Yќ%Di�B��~T|�-�4r"��*��h�)�^�Q8Z�Jr���Q�6�@N��<�ǁé$>~�7��X5p��[�'f�5HeC����5I7E�U-����&��܄T��6�q�6B*;%:�o�O�x0����EÍ��ݞ�i�󺯱��T#&Ǽ�e��ඈ�)���K�H���r	�&d1xQO7���-�fH�+yͶ.�ͿcM�O9a�9L&T&��r� *:�Ձp�
�%�Dܲ�a����dh��������D5J��l��6lQ��IZ,N��F�~�FJ��]��_A-@�Rno��_=M��F�he�T��2�H�(?qi�Ɉr�ɜ���ѧ�'�7�X�!�\P��/�:�'�-��٫ޙf�+F�*��"��(B�C�Zy �\m�l��Sf��HyA!C�#�
�v�P�� �B{�������gEv���V�.vN���ێ頍�r*�-����܈{����
o�{��$�x�d��0����2? �K�&����ZU���)�_A���x�:+��Q�
� 32�'�Ҭ5��aAꎷ��d�6�?@+�����/��!3H}MK��s��RI�$U����W�"�9�S[�u�~yR� �n��ϭ��$���d��M�_��e8�Ÿ����!w�x����s�q�@���#%�x�q���ӗ,��րH�2,���-8��Rۃ��6��v��M+s�ڰq��f>����"���d�&6�B�@g�3l^�����G����ATf�7��V�#�e�'8��j �r�7V��L<L�uJ���J�h$"h���c?!��)����6��Z A��W�8G;ꋐ��f�`�򂑗���M�Y/*�ӷ�F����@������,���L�2�M?��8n�v��W'����� �7��:��f�)�j�*|��gi�3���7s��S�;��ܷS�����3��*�ʷ�A����v���Rad$��^'����BE��Hi\'��ZR��M�]N��y�H5Ȟ>?!-��.��i;�w�PC�9�����}���Hh��{�T���~QxVf^������"Բ����ʖp!Z�����/a�_ןEV��  r	�]��}��aQ	G+,/��쵢9�z��{��h��rI�>E�m#F%5ts.uuYE��]��D�@�pp����3��.�:�n�i�X�7���/Yn+��_:���X����-t}s+n����u-��9�!�
0q�돣S˗:m����О������M5 O.�^�*-K��9Ք��'��IդU�ZƼ�!S�S3�^ȷf�x*�*�^o�@��&&��m�s�sPYD ��ol��p!"�Hr$���w���U�*�7��_��$�m���~��Vh,Ù�2�����jzE�� e��9;��G�S������~�Mۓ�)��:oӿ��ѣ��I�8��>��3��o�NR�H !]�1R��;<�b{IU�p��4`�(��J-��[ĞM�TCQ�T�xi����"���r�)e��7��vDP��q(�#�ʺ�H��͈����F��_��uQz�&v�-����7�|�j�켳O�&����A[[�x����ss�V8K8�i�%�A�?e�ڹOj���Io�Wr��9IT�==٫�0�L]D��q���Րn����[�Y���V�(��w@�Gy�OEP�k~q���2ᅭ��a�Z��:��Uc��P��%��cd�!���xOZ��=^翍v`�[ȵ�ks�ɒ�yܲ�>P&f�'b��e<���ߓ"�����J�f-By�A=�h��$��}3\���AH��S/P�_48������%�����j��?�P�?���C��h(h���2�)��U�w���,�K�:7k-�-��:^o@"X-��ϝ�����|� ƶ,�M����!UE�+�=\��mt��|�|9�c2�X7���ԟ��qhG�-W�a#%I����tDwﲡ�0JP�� �2|��T��hF!Ge �o�Ͷ��It�e��LMMi����E��jY�=/��>�QÇR~E"�N�UU��G��!��Z� ��%b��kbT���#��tU�I:������P��$S���>8����4��J�cY�M|�i[�,�z��%~"����a��<��I����=g�ep�|!q��G��-?�y�m����xWX�R6����4k��wf�u���K%Mc�e��*z���Q<䕠v�J ���I���D}}��������O��KG/���R�-�Y��M�Ѩ��g��e5�Nm�Km��%�ԋ|C_��r>e��Y��0ڙ:�;�*���@��l^!ߤ��v�6A�z�z��牠�W��^��T��St[֤�C8�:�a�O��V�0�i�X���Inz���8�2�}A��0<�X�?@��p�Rwy���3�
By����Q�	�S��̡EW�d+A�}�QG����;�IX�f��^Ʉտ$�"P������Q����E�d�̍jC)Me��L�0�bi(� �(eu&�͞vQC�y�)

�vgT"<�g�y����<W�%���:�]�*�9>�r�/Z,Ձ�����r���7n4H1�F�cR�S��r��7�ـ���������3��俘��7uɐ�?e��g�!]X:@@�ǫ+�L���\Ẳ�� �y������o��^qWWk y��
�|Rnj����_3����%��#.��r��(�H����R�VǗא 4����^���XlxVHYEB      e7      a0ч� 8#�S~q⾺����~BȴU�ƙ�I����Ӵ���Q�E��8.K�mtv(����m�?`��t�IViIk��`h7�r��.��wN�� ͇q��\�?��EW�������&;G����F���k0F+�D���Kd�����f�}:r�2