XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��@�y�"h0N|R�)�i�!�)�ந�AJ����hfz ,h-��j��/rU�n�"S����L(�}�G���]F�F
�Lk;'ړSJrt~�,�D����<����}ص�8���.�n�ĿV���5h"����2�����)��@>ئI(��$����܊� ��M���<���[;0A*'�-�j�.�Y=�TtF�
Tcz?�>��]YY��~u�1/?g�{��J]���2��F��J9�%hMRZLϏȟ�M����-��-؀p>�,�),�L�2l	�*E����f�ΉF3y��,ڛ�'�����\W`ʚ�P�X�$�f
���#�X,�zU��n��7�Q+/d.��Ŭf�y+�_l\E�e�+�Z=�N�f�F�h�1��|Q&��/Vɥۃ��v�-�
Y�V���^��r=�-�}��}��r�4�	��)��L���?!���67Zhim��7�1�mY�}ʜ����̅IZ���"�/ۜ��eW�@���}���!�3��mU���D���e�A���-LN7���>�0�����#�1$�w)������M�)c.�}ژ����>8��K������b��7�=Kw�L�����uoN����8���t��=����ߥc5.���N��_����X�A|%Qy�ո��QB���u���=�
�C���b[���TgT_Z�]+L5��QF�gm�ˊ�����kγ�<�$B���N�mj���E.C���S};��+��c�XlxVHYEB    fa00    1950�ո���O���P�Uy����V��ZJc��+�Ŗ�(��b���k	
��y�Wy�3��҅� D�h�$	���M	�ن����B���������V�t��]� �-�1�L�T�<��_�Hx�DA�W�S���6�;ċ̎����41��0/Z:ʁ���S�WZV��K��%+�&T*p�>L�'`5A)p��E�����@twٹØ��f�Å���oqh�wKD)8O����0��켵:� �6�Z=>Zz����t����(2�/�x�mҁ�q�bN�/��bn��ê�`�րY��"qA Y�
ۻV���G�(�/	�F��+8|~��'wt���T7_���w���xa�:�^� 	цr�.(ġ��;B���DO�Bt¸�܈[?���>��;�P��0��k��
�'ZC����y�K�(P�g�U���BX��ze)k������k�?���6�<��W���8f�vm�XZ��_�g4E-{Զ�$	�����*����ê�IFz��'*'�oYB�k�+�Ց٘Z���
�o��S���,�b���� �^�j �Laԁ�U(�8W�/=�煠M�c��@�=�$s�#<C��v���,�r�����Ny<��~#����Q�A�B�1?%���FN�1����}{��;8ыy:�MϽ��o��']dkQ�h,tx'O���04 ���]�d9�����zr��\��H���}"��h$�������~�K�;.΂��~8��-�m����07=0M)*���z?���1~+�N?<Ջt������6a�W/�k�tB��a���hw�Y�1�A
��NpR� �G���8�ӌiL��8
~	,[)�"�[X����uH��xC�٩6o��/��$^��5�`���t�[;�ͻ��.���|�`h��U�"֣�A&�ovˏ|�~�)��hS����8Syl|�,�kE��#�� 1�zL���Ɣ���f�|V�O��'���!4�tD0�xB����&��:��T;l'5�FDUZe$�߼P�h;�� �K�T�=j��qI>����
%5D��aRZ!����x�} TE9��/1�k�C�7(xv&����cy4�]����y�|��w�*�?�?����m:Wy�s3����������P7��;#q4=[�L'�W:.�P�������a��;[.{?�2�u�'=���a!���.�d�zּ�q5j��� ��x�k���������o���$�nрŇv�6	jv�Y�i!C��!���*�l�l~�Q&6��ëB�r�1��h�ᴮ4��*�V�VV�I��k"�F|����&�w���Wi����N3~��@�=Z�ux���0I���(���Y��HV:EuZ�[�j�q0�{�V�~�	���a��V�zڕz.�/[�<�/�Y��aNp_`�%�I�M��!{luXb(g���@�s�k��_\iF$_�L!ǜ�X��5`Dx�/���3�(��&1�E������oI�p؞}I7Љ���*��Z��4�r�c�.������#���]�2$x�n���.>ȿ�&N+��`�c:��}��hq)����sZ���1�{&\�F�\��jE�y[��p�*.�؂SK1���M뻎f�s-9y���"�]q<i�0��}I�
�ue7u�`]����	�8w����~����F yn.4
b���(�S��M]�����$�&�s��%����aWvQ���^U/ȥhs�B�����
Ѱ����XT]���T j��/�jiX9S��ʫ�y����Ip� t�1��i�W�3�����4XOp�� �q�tw��?[Z�[Ŕ}\[��Il_T�Mh��g��&�m�>���2��!�U�����^c9`,q��o]Ԫw#/�����ic~]��Cha��8���q�5�i������?0j�l�r��s�XȰ��]�퐣�����A�!L:�9�x��=B��:M ��^�V�!B�W;P�� l�>��qB�F�)i�V��M"�ZX"���m/�=��'`�5-�-���3�.1����y1^�շu���(��MwSXE���leT��e�n�_�;I��7A�.aj+
_FQB ]S�Gl�T��;z�`3aa�y�a���0��r��N��z�.AK$Upv'q=/s3��;O�*֋�p�钞O�SX���c��	|�y^Z�Hދ�H��<��d%��v���7�ރ�1N��U� Sܵ���ϸ�yg(�"ѝ �9N��Y�3��}��I���0SԮ�?7��6amI���	�dz�_�G��L�VT���R"zr
�r��Ҳqp��p1��K�uO��bf�;�k�7��߈4c�}RC�p����z��"�Of~2TXB>E�����0�)�S�u�@`���؄U�:5� 8$WT�%oЈ}L�������Eem������J�B&"���&�Y�D�AŵG�g<_P�Z����e"�|�N2�|��s+��2�ջ�D7�ċ����!�?a?5�3?
��Y��
�q�!���Vs�7s+��.&�pC;d���%�H�fE�&���f��i���9�ح窌�<,��rLej�_ �Z�BU�j���V�P7�`�����/?�	�-C��!l<R�?�6�}p?�v��|h����c��QN��(쾷
M�6 ���;�6�D=�çh��N̓O�ЇW��F,�8�!E	F:dz�� �&ɤ�6D�$� �痣�d ۇ�o ���a��$�r���4^䚎�O��
����)����Opń���J[�I��n�R?�a�E��˖�@��+wL�B�������Oy@w"a$��0K"��⥘���ĕ0N�����(�S�,�r�9�9-�o�ؠ�;$��22ӑ�����G%c��'��,��+g9�$�6�c�3�5���$�5jzc�v
���otJAk5&7���e���0�Ԝ�������A�Zp��fܨ�鴥�/�GU<�o���.m�}m���ͳ��Pd�G��@'�9}���u�8�����[G�K؇:Ȥ�0���;V��� ���W�oj�s���?��WKh�TފD�.P�.]#��6[�U>�ĦuM�/21 R���N��=��r�U�c�*�,����h�F1.�狘�Пz�-�ĀUp��-1���TR��۹�0�ms!�;��jz�n�L�E݄<���LMӗr��R�Lȑ�O���X#���^���&��cz46F��C�v��$���5E~'�KSfz��I����T��.�C"���ڰMO���*�4S���0�ãw%�m ����>4ug"���_~]f8����>����w�rI�As���:��O1W
5>�7++h{�U�œ�S�>�� ��	j����<�Z���-�uD��xJ�_�CC���;{���3��&_�i�A�:J�:��!&𙂑�Ea�����[q?Ģ����b+g�iYO��2��������"�u�k\Ǐ�F����h8W����5q&��4�`L�^XTׯ,(鷧/�b(.�N��"��������&���D�Ճ�u�x�=�5�[F�-D#Ѐ�;���g��杋�b�(]���Ba�,�}[qĮ�ec'��x=7 �O�~�U���zgp���撽C����r ���1��D�\F�dB�
R!�f=���k:c�R��� ��9K�k��U�w8�����G�6Q�
��o��R�?=L��OQ���M>*�m�z���������K���Ų�ipR��|�)U���.�-�-�	S��&;�H���e����A}kjJ�}���
����Br҄H��<�����zQ�r�G�-�^U���M6���z���@t��skq�R��'�3 Nڝ d#\��[����+�IVu�����e��t5Se!vs|�`S���3h)��:�+��sۮ���:�`YwR�LY���q{c����	�ǐ@��=�d��EY���\�d o:m���3	&Jچ&���"����?��f�P���cٌ,�x�*�n�а(]T���^N]u�q2H�M����_�~��
���L���dr�#�
,ʡg����3;��ۧ 5Zi����ˌ5p���T�8�� 6��"�'����^���X�D��a���F�rYܽ�Μ���E3��X�Ur�O��*�(��M�NK�:�ӁP���"��c5�uK�/ B°q�^G�-(�)t\ Lh�`sOX�q�b�-�p��g��(��.8���^2�Ԟ���r�
�VU�-�*.Z��U;�?K�՟ES��u�"C��47[�x�����������}�0�,?�}י�i��������S��5����.=����e�u(�o@�Z�\d���%t#��.�JYS"�X����c�vk�`�qN6�o��V`�DЦ�|Sv�Y��1���[S:cK�3 ���!	o.���o�cdL�sG�_�W�:~W]���K���}���N�[2��Ǭ��gq� Wk�fA��=5b���� z���h�&�OԠ��X���Q����@u�K���:��˞.�28--�i �\���ysq
v	
eD��6���O|�[4/��Bſ�x3��Z����(2_���.��I��3���Uᢸ̗��q0q�ÄS_qgYY��qd
E�бfK��F��Zt�R�A^�J �����=F�J�8���ǜ�Za�e�]L�	G��'/ۘ�K�5�A~�B��!��̃�JWQC��Ǧјz���һI��u�)�
�^�����tYÁ%��5Nh/P�^�)��ǝC�dwy��MYg6���r��TzJan ���q�	G%��M��w3R�*��g���Ŏ�����H���h҇أ��7�u�y��Ⱅ���~ɋg8îxF�Plנd�uc�Ң�ll�Ά��i���$}Y��ѩ��ƃո���h�����&{A�-o!�wݵ��C�h�m%�����-�k�~+>mM�;��oo]��	7�I�x	��y)��}�'����%���^w$yUB�al�%�8��V�Vr�(C��0N�#��t��f8dNΚy�
�ibօ�A${�5	���wY�U�k��j��5WQ��N�)���V*�O�QV �3k.2�R�&9x����LӍ�?�P	o�{�_L�#�uYh�j��16���h�"L�y5s��~���|U�?�q5���j�������< ���b;C�i@���$���Og��wB3k[�a��D]����])�@;�G�9�B����R�2��t��o�hѱ�8DG��n�?�Ki�,V2�S�:�- �W\�\X_�9吐�	���<�a�H͈%��\!�]��; O[�����2݄^�-�@Y6&
�WV�Z��c�T��֌���%��L�U!+�7v�O�5N�Fh<jM��t6hOٚ��P�{��i�'�Ð��� b�~��CJ�����쓆������T�/d5n>����u��H#�[��;B|;�邜6�k!0@��nø�54t,��v %���E��Xx�4�jE�@�k�#�������Zz؉� ��u�l�%g�����o����/Dj�4�%f�w��dA��e�K��gb6p�|Wَ �T�4�KXh�:+aD,EuKXG��Z��SW�38H���u��3�Q/@�v�<3���(�9�����`���� �u`�������F��7�b�H)wU[6*���uK�yt�Lu�:|1Q��p��PbLt<�UУ�<[�a[ �r�m��h '+���l4j��HOS�}����m�� '��h��ʁ���N����tԫ}D�;
F��T��a���OP�
4�3��+��Em�=�L��蟣�-�O��e�S�&�0v� ��aC ^l݌���cN:��,g�^iI��3��s睽�4�Je=ԗ��������g�	��!Zl��Au"1F{�"�GRY�J����Cc"�WS���~W>Bx�T!���@������e�e}PP&d�H�������͜Zw��+{��^�������?���lD닚S���"h�Ai����fDgVh�tQ��c6�"���:8�(�d�E���5�L!%ű�ڕ�
*o�!�#C�B�p��ņ5t�Ti����:��#4��)��`8�%4�kX,5˙U"A�<��F=i5<�CX�b���}2��(�+ �`I��%ߧ��U �<̩r�=��@�/V,ψ6��z!��=*��tU;��@
�L�W���g�&�򍛇 �Ak!���gre�����`ΐ��l@g �j@^%��5�����:!?w�<��2/x�Z�`v���CNRW`�:� 3c��kr�Rߒe8Lz��7�j���/,�[�Δ���Mz�س^n].
�F�L����R�؎�,�_EI��6��`����C2������=c4�vJXlxVHYEB    fa00     700n2ظ��\aA!d~.k'ræ��eS��W�U'�	�Oͱ4� VrUTd�-�M<���A�
��t;����T�ZB�Y��S����)x"�7�5���T}� �I;f�N~��@�>w��lCQ�qHXΡҿ��6R_���:[���b�����QW[��AP��I]A�?�x�D�&�$c'|���8����D�rI"��.��� ���;/�� �e9z��0�${�(�rN�a�բ�yꕨ��2Z	���h�ǇM"�Q|���XM���$277�����WK�E��Rt���h��FB����bgT��
�0]X���2���苾�
�0̎��	�BI����	��@��)\ŉ�3���}ofk�,Z>���i��\�B�`��5�����0w"�-:� ]r�\�u�i�>az˙�,a�R�\��'���=\�,Ga?K�61�@+�J;W�G�UL�D��`����PR{������`\�Ȗ�pѥ=��,�
��Y��#'��^�0~��ie�}�~��4нhK���D�M��Ӗ�J]���ƹ�:��4� �aA��E�;t����Kj�3=mۆ{()�$�:E�23�G������K��VuY؊�2�A)��-y
���̞����l|_����NdP%��p�N��m�yKh�@r�둬X�	��
��(� N�8E��=��\��뭼���Fi�(�t��:i2I�~�F���-�	��/鞊~ө�w�V.��,Y�����&q�s��c@A��_��2}��L�v�Ϡ��!�-c��GH�R#�8�����X�h�,��*7��_L�;�� �o��5�.M3�m@����e�aA�8Ί��El`� � Y'WRId��L���[�W5b���'�Tڛ\�i��)���ñm��0�Y�X8�,<��/�M���#o�|؝àu�IXy�?k]��)bb1p����j��Q����1@��J��S�Ux�6�T'b�ך?�i�,��E�N����叧܌�ֈ���9��j��*�����q�5�6��Ė��9��e��L�Am{Q�����O.��� ����|
|u�1�V�n`zi��|Bziz���J��)H^��x�t32�^�hF%�/"'���~R�晘6��Q����۶�=�v0&�Ah�.��RQ��2����g�����������?#��QmT�~p�w����w/6�G��;��l�@ʭ�]�^Qe�r��b(�Sq*y��K��UA�Q�Y�ݠ.�����xD��4��%n��#��O��W�fxb0�`���e���Ͽ(&���� W'���O8����ͳ�M�p$ܫ���A���� ����d�$�\��� }aA-��Yg�Qt0��+�����"�o]�=���d��jھ$f6� D�����/�#�+���!�T"#3�,,��"�!���Td�����s1�S7�8�����$��\T4h�)S�����5}�1��D.�ׁ�	)����d〔 �ǲKam>�<��H�.��;���� �GVd�\��.Y��(Z:�Jz�w=�!��&��Y�Z	�v����������e.?Tꐂ��Ai(d
�Cb��z�Vo<P(mt��%W`>M�b�Wy��$��@F뛰��J3[q���Y�#&E�*aӼ$=`�7B����Z�Ż���W�X���j�������}]�A���<xF�G��͌�{�Ȍ�ɡ�"!Y�M6�����%��^�<V�!@�'eֺ��KUw��"p޷$d)���W���4:�q��#/�g����TXlxVHYEB    77da     a60�n:�R)��׾&<%8��8�9���}W_H[c��e⺐Br�Ιօ���]X �
:EG�c����=�V_֟f�~�H	ښ��b������ܫ"̪ ��� ����K�j,�
�p�$���O�l秪ۍ;Jۻ��_�8��n`�<��&\ɐ׫� �Ы�������O���������U���i\�Pf2��JE	����g��u=N�|k������7�޿^-g1x_
gt������X�D��At��%iɁ)��(��Ft�����`j���ʼ�pBi	.ﳲm�T�{1��P�g _�27��LcG�h:�v9�b�Z���rZΓ47���(YD�v���q�U_�~����������I�C�X_!9ɼ��	*�ˇ��m��2B� �G"8��{������gχ��a���Sh�jLEs{%LE�p�ś�5�����?���Cld��>��.�\����4�,ea#�$:V*>����`M&�^U��z+�L}�Iy�����^�J*�2���'�dt@f��&vΚg/�TB�+6Wza���v�s��~S�`b6��� �K�]R�`���x0M��ѷ}��@l����"������+^+���1�������^5;/�%^��I<�Ȓ8B+���X��8�J��&���(�/J���N�Pm7�Hk��^2����3q���F��F'��8M�dY��W�tX�O}�[�CH�b �G�թ�d8� ;�tq%�!2���4�ƃ�*L�/6�+����P��<(�*�Y�-��u���y����-;b
�����eֱ�����+_��?����������O0s�����o *�%-�ӻmn��^-�c�NP������h�ē��-��~�r
�;C6��|�R��qgS���k0���\��b��%���SM��'+���$�J��#������/V�eS%��YЖ�:@>�&��T��z 8ϝ�N�CI1�P���� �f<��K�䦅����YU��vD��X��5j��W�_��"G;3{&@2n~��-���1�����'���r�k{�bgs�\��U��ZD�$�h��i�_�o�s���W�7��If���
*\B��	.�Y��>� =�ǂ%)!���Ͽz&ߍS@������>a��m����I��r��:�A���������ԅ���;��DZ��Ld�fd��/Mzd��f�â���rxB��F����CៀB�7�q�o�Z#*?�Pl�;��MxB���\?˝�À������O�U�o���&I�@���e���������=?|3��i�?�{�]�iWKx�n�7�ë�tY+2
�t��#�lU�m��%�c���s16�YIPwd=f�x��5��[ ��D���p�Z��m�'��a�^� �iu���`������Sh.�-�g
#}?�z/�OY~1�^�	��v��,��i���[���K0>�!�R|e螡]����I��ց?G:^>�(l9uô�T�|��y��A���x�ٶ���kXT���a&�Nz�-�jE�q�P�ϱ�@<c�s�����[%6�#�L�F�ʦ�l��G�@\!�B^p�+�*�b����R��sO5�s�Ҏ9P>�y�c�S���LA-��i{'���Ҙ��cl��9�{V��~�Pp_~ST�٫�X��{��i8��Q�\�u�����p�H��&�(g���@#�J��w�[\L�u�[����:�)�^�r�N��hR=(��T�Y��j ��J�Q�-���#qg�:���!q��p�/U5j���o.�)o�꿤Y�R�$�c�~5���y�񁲱�]��V&+tҵ6 >]⭠�v@�; �9��O�+�͂�ȋ���!%��I�rn���+��W^�I�M�m.��V�o��_�ƮD���}�>�����\F#�-ܕ�Ya>��R�_z���1pR��No��':n�#�Àuߍ���-�A�=�����������c4������(��"rଭeQ7<-_�)qN���i5j�3��U�M�'�S�^�o�|�)L��뫦ʿ�������3��Y����$
��|[5��n�Y�壓�pE�F�R%��#�Z�d�D=O{�  �,ǋx��~�c|�_z���CUT,
���~j�I��`�Vhc����8�EdP�3�v/i�����f���[�]꾉�#B��a'7�L�ēѭ&͗�	��=�_}�p#��[��2��l$����/\*.p�X�����}������ݡ��0��_��Ha
��a����B�/]9��z��Y�5On^8o��W	�Ӏf��o_ p�u��0g�g��[�VuARt�k)Ɠ�PKTb]��v��܄8y�A�K�p�E�����ΙXm{RR��@�"/�U#|�%��X��t�xv]PT��}�b`W��Kp���#VВCJHr)� T{Q��jhR��-+[ew��I�I~�_��W����0�]=����n�7��E�p��o	Ҟ:S����-t��;-�\����K �ɱ(H>B5��̎��SE�C�A,��0J<��{f�h^���>�؜}
8ffV�\z�Is8u���
��7j�PA嚜`�%���a_ޒ�g��bp�v���