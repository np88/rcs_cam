XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��5Q(V�����cy�ʺ86y,LNU����F`u�z{�y�bg,w�� ��q_��؛��N��>�[t�{$5[�۝���p-��ld˾����G�K��,�em}�X�3yi� ���Zn�n����3E�����D�u��G�}��]Yٻ�D�@���N,Qk�b�2�J�'ϛ���i�dF�2����V��Ϻ�Xr��t���F�J�z/į��J	��c0�B�naו
�%k�g�"�f��l�1#t1���5��/c�t8�3M��)���H�x� �����ruP#b�9�;'�\��?w�Q л��kr��%���jH����D�U����6��h�&�&,���t1�h����6�5���7ϻ*}9��3U< p;�ˀͬ��:!�D�A:���.�ݶ�'��k=�����J� ��K�Vߝ"v8C���]�?o9���G��:�U�Qd�L\�L����b��W�$#��hwu���S�|Gߘ��p��{�'ZiQ����Cr�RP���̧Š��sb��a��1��Ē�0ްBSSa�u�\�R�� ���6���#�#j
_��ƒ� f�.Y��/N��a�M�jHC�
ߕ:։?֛��CC�X%�O�:����}��i�j��O+aN�#j�Y�ˑ�x! �z��:�ؕ��O�çEBB��UΒ�Qt ���.�.�MwM�Bz+�\TG���T�~;�0���2k?9�p�,O�����hN��K������!����M��~���nŖÏ�?F7K���XlxVHYEB    c6d9    25d09�1��=�3L�[�-��@y�B��z�0l/���E���l��*�x�k���+����
@ߥsd}��X{�@c�1gV�=�4
;`X`�+��޶mu��h���/CB"S���c��4���N��4B1R���J�Mo<�SUs<�G>i&&����`)S)j��&R���@�ٓ���]����8��6�L�q��W�S4�n-i��i���	��ц�zA�J���d�#8K(�����0B�^�����%��Y�X/��x��g�k�!��it�%c."*'��z|��U��IB��cJ��n�R�7�A����܋��t]��'+Ӊ��m�r�DG� γпfO��h�'i7Eڕ���ټҞ�}(2�gy	�:&��-���k��z.��l؋{��� ��n�}�2B�ʩU`r��������O7>��Go�iX�D�ċ��\y�oUa�mG��V�*6lV�ŝ羼"�f��1p�wVݤ� �N�b{͙��l���aY�hEKٮ�9�k��0����Y�ԡc<A�,�l������DA[5Ú�)cRۻ6&V��ӑ��c��Sč�of{Ğ�N;�`�j��������3;�����U�J�ބ��S��?��L� C�o�Td�^sN	��[(#���c����Vt����e��v�Ve���l�?F�O�sd8�bSr����,�a�Jѥl=�/�M]�5�JՃ�Jcj�3c��sZXdδ��Ǹ0��G�D��|���R�c�R<a`[=��eIҚ]9@ɂ�w�4�L���P�s�Nh�S��7����� �8�݇+p]��#.����wUޢ�J1r,혧�(2��p.}����b�0b@`
��X����PȟY��\B�J�)�}¬��Δ"�����������O���:A�c嬁�+}��z�G֢Dī���Em�κ�vEsm%�(c������m���Z�P�c:p�+���ly�����wND30&1��<��:����Z26هB3���ع�Pi��&��+�v4���$���@�/�C�T���\4�m�GA'0-��cY�f�u݆�8`m<7�o��v��:�(Y�8	�ڂ)!m��]7{����F�>*h 0d��<���ؠe��2(�M���,jm�@��B|�"2V�)(�jR��N^�����k��X��M��50q�h�����*j��e�}NS���7)�Spt�{O��K0�קfѶN|�H RW��ԥ-_�K/�Ʌ�����V��Qy�g�\Tf���e��<_=w�����Cμ���V:�67��CD�J�+�e�@��AK`�'H�1ɔ������Hhed�n-�`NԺG�ͻ3��~�tœ����l)�ё׶4��� �M5F(�+�.B��Qb�כ	��К�Y�8&�8B��Ơ1��p	�F�O�"0���U��:���s���iȠ�!��|j�o�x��5�������/o_�	`��!ϝl_��8���,��3c�i��=�,&�LԻ�֘���3�M�$�X��\R�l�5�s��r�ET&�s��Ы���"�gSN���+��Wk��_������%�X�w����X����-}a�rk2������|�	�厡��vgM���1�q.t��!�쭶�h��:��t/̇W�)F[����0�Vo<c�\#����4|{�+�M�̕�Q�\e��6_�%(�: �H%��l58�J�
I���l�Ob9t�F��T���X���ǐ��D��K�aU��GW������{i�I�Vȉ�W.uA�dZ���;_��I���ӱ4?�|�����.�N0羦ߦ˩0M�&1�Lv�"��u��~A/�8�A@S�d��õ Q�8�T-a��6[�D�,3g��E<����Nu�6��oÙC�4�tt��NgӷW��0��8X'Ѣ��jheC*�X���r^�I؂u8a8m͇�µi��>c���a�j�52�餥S�+�����]#�|U�!8�UbM
��HH��'
?����z�������=��J�`x�f(g'�3(��@=	s���qd��cʌ���[���v��t���V���r��~py'�kL��D
��f
���`]^�԰�D�a��W80V��/��R�`�2��#,��;M=�m
9�|� ?Fþ,��_��!3�͊�[�!wѺ��y�6���r[`p�.$.�w9�'�Yo����aA����ʞo	�Frτ�����'K*�p�?�/zN֥�����5�N_�b`u��}=L��L�IE�=��n>�����'X1�Yn�|�u�~*��K	R8�^\
�euCa#��ԓeCF��Kf|�C<�5��q6��9~P�4o���H:�W���}+ꇷ!�,"���T�����#G{��8�����`7�c!o�	�v"��q�U���r�r��O��_H�ݰ��CP�-��esa��L�C�ZF������<آZ���[�oq��C�8JJ���X(���@�E1T��{�Ds,��ݔ�W:�حC�_9R��wBM�l�k�3���WP���Sc�ں��B%�f��Ӭ	﫼�
�bѥk�4qs��_j�F9�ޗ�_�j��bTe�/k��n�-U��\����!:|���ݮc�5�]��7�
�W!}�g)pk?R�%$��l~�w�����x���?���fJ>�g`qMeK�,mfeBwڔ��v5�:6�ǾX��n)n��d�� 1��Y����Rΐ��s�8���?g�S�L饠����Tf�.�u�"�|�?>{�|⠳�S,q��+_�NԂ{��vvD��U�q��E���ZqbY��X�<�M�Y�Ja7k<��i&�k��e����o��D�����Wș!�σ��܉�����n��ƺǞ{k�3��#C����>�Hf���o�,���|j��u���^^��y٧N,�c0E���v� �G�Z�������E���Dz���#"�z�y�����\E/��SX��~Ɔ��v6k9���;�ۿ�ށU�eߍ4�ѮqA��Ά@ZYf%X��G]���{I���?bcK2Jԛ�����.J7�h2e�6��W`x0v�X�t~������>*�Q3n��>�U��p�J1��z�V���r��]eU��K�LbZ�y�c>�W��:�w ��1;n�o�*p��MEʳ5E�J7`H�G�g�p��=O̕4����>���I1~rv�wCS�}d!0P@�a��~����>�z�'Bg�
Z�22|f���N(pp���]�e?�o�x����r-�)]	���ً費i��ҩ0�����/I'hSu7�+���ډ:�"%�O�q6�!��'�� �R���8�c� ��5�g)�3�`��@%_Z�i/���|���&虗����rX�a6	ur yׂ�~���T6w����H:z��A؈�a��p�8�{�ۋ�?�� /�e]��j��/p8�܈-<?s�CP��X;L�5���}dK<�3���X��X����Z�6ިAak�H�|�6�`%?8/�T�h�	�ٌ��a`�%�n�����g��U5�j�lc�_��v���B��D#��ك
j-([3R�X�R�+5�Ht��a��x�tVW�R���y�L�>{N��AT����C�e�F�����-�(�#i3��vͱ<{��H���fۍZ�ͫ(��<�v"Bǭ��J�ث��*�xXs[��Yj�J�&]Q�{�i��x���3����oP���\��6P��)����A1�_�p�!���'C!�B�CB�z89�{�T@�ɤ��	s�V�7p�ʽM��07����n�U�?X�þ!TO}����*I�k5PU�,I��/��\����i�<4�?N_��7��9�WU$8N�\�ϓ�g�)i�
��S�Qoq���5c�k(��%V�Ǐ�S�2��d�W����^�4I{���.��L]����>9�Ԥ���`��)֮�v�z�ݹ���yQ��ym.����Zq�M��*�_1�.��Q��;���YL���Z����xϚex�g6X�����V�s�TO����|̠iɻK�Pb�ҫm����e)Ta&��4�?���AD3�-U��%�>�u��oP�;�!�i^_�6�o�F��������qԗ�����fƠ��Y'�\Ϲ��T���=Z���iS:E�=�w��e)�?�*���6����a��cg-�߳FE�> \��~����۫���|?��V�Px�S�$��V&���X�QljK�U	A�xL��IJ��{��+i�-A\��fY�
���;�4�Ƃ��s�t�68�����Lw�A,�d5ub0wijҋ����ܜm�E #�~/䰍����O�ǲ��6m�~��\I87>IMV'�/Ƣu�4g��YfF�8�S�"�>�����?^�Zfz�t� k�n��%h����Ġ�(���}z���Ӆ�װ;~�#T8���1*������C�h���	��L�W+��;�p��zlK]�3p--��+F8VX+�7=���<�5�⨻t�OY>�`FRuG;Է%Փ&�FӬ��B�_�0���O�(ym�|r�U(�R�_܏1����u����\>�Cw��yJE��mn��X�&�E{�����Yry��'{��VL�+�U@kj��k��R{�� ����5�P<�҃�54/���/@�vu1 Y���&xKT+�z��{D���R/���Γ�6�֠Am�����:��ڧ]5��}	+zv�AJ��@z;�_��ʶ���y�xm�G0�z:�D�H�������N��-��iR�ZJ�&�����Չ/����<Y�Cs�=(^�Ƈ��{��t����T6� �
�bM��w-l�Mp+e��Y���PN���eL*�] 0�}z�b<�<�#���'w=-N�_C�dl����O�!/(ͅ�C M&�[�r�E�������$�Lmv^x�@���{�_��㱐�"�п��}�Tm`��äl5�1ɝ
÷������k@.ً�Td�wbb&�a���-��lP�Ҫ��{�t��*of�XA ���5㠜��
�"��> hw����QO����n`�.� �}�T�p_ښ7�.=���}� P����L<p�}�%����_���O�P�V�}[  +Oc����~���G�B�K�D:6g&�f��5�,Gq�N�Ѡr��؎�+��+J�,�M��si@����ZS�7�� ���+A��p�J�a>!�<m���fiJ��J��.㔠E:�T�3��sɌ�}\3=6ץ�R���	��4*�v/`�o_~%Y�j�j?�U�A�&������-�X����u����N��F�³����s�}����u�gE8�����ls��\ du@�R�bt��6��#�R��Kbq�'Fʨ��U�9��	�A��m�=��2��",W���+? �����ݵ�=�3�8領����n������c���Gv�T4=���m3��6�N�W$��L(�S�Ό���e���J�� �V
�.��^���v�Lj��Y�y�|-�LH%MQct�X4�p�Nbe"�$���²���;ԨpR}�s��.��==��7h�� ������+�d�n:�v�N�fuE�G/�[���3hq��~�1YF	Dm�x�v�H�s��f޶*��w!�'ڱ��Da����}��M,C�x�X ��=��g)��ܻ�L�����bD��\��6����`���D/�N����ija�9Hq�&&�Z}!�݋[�rD$d�*9���K↟�Z�f���<R.6פ:�����/ ����k�2[�ia��A�7&0('��<�x:���xNؙ����zΉt@�yR��ϧ�s����/���+��9<(��w�#���I��G���*l^��p��kBi�P&ћ@���j�$��fĝ�>��a��(�xH�OY�R��	?H(��Ⱎ��\��.��DC�}R�iO*��Q�����,�`���Uaޘ�]�0�3e���8_y�Z�bx'V��l]�[R�q�ޑȬ��Zk�P�^�/�
ׁN�Y��T��U�d���N>YZ0v3m9��d��\#��Q+�j������I!�ZN@�)#�j����-���D��8'8�8��g�uFg$T��6��j!�'�i�����⋹�DZ���
���w�T��8�Ԟ���$�P�E	�XD�k�$�"��;�ؕ��֪�*��0�Jf��;�у \��_�ϝ�T�-��6��-̞g������ü����ly�̌��AN��Xz��K'[�n��K��f�ދS:�l#�;��?�P1�ݜ�����/kD�����������^���� (��^W�Y8������;}�_�h��<Y�Ӯ1Yo8�`��ʏ=:{.Έ6>��>\+K�(�v��Q8�F�3��~�E�0�m�ש��V�W�#u���Ma���`���tԡ�88͗d����)�uP!j2����W��~��S�7����YcQ`���z�'z�$3��p�{��v�8������0	D�_���pl��.� �Br���	H_���W�%V$�KK��������u��	��/��u���W�F�:����b92����(�xp��	�蓲|���ƛڃ�Ʊ9��6l��l��چdj��R�(��Y��J��i)n[K���i��C�]A�[4�n/58F�Pl�Rb��V���[=���?�I�~�Y��R�*�2��V�Yx�SJӲ_mvu��\�Q�|8hs0��;q.$~�`�@�BG���T1�I�Y������GL3w,M]gT	�/��1e@p��i�3��w���<{�<xM�U���Xz����D��oW"*������߲S�'SI��E;�x�=��4\�sC��.��b�ϥ��[73qG�nW/x �`v���U��4̱�Wx�䖅�{�~U�4�Գ'��)�x ߽9=;�g�a�����{������d��/�WR�z�
�)��DMo���}V����,wL�N�u�_@"tt`2��L�hy�hp�ȑ�>�xd��:��(i�/��'*�PH'�~�C�l��:��ɬ~KZ�'<
5�Pj\!}'k.,+,�J6t��!�γ� .�v��p�}�:����v2��4��Qw���<-+n�sq��<��\�s<U�!�Z�3�zy��򯬸��p2 �&Uf��-�/����4
k	���	<�wy��6�2S���kU���$!���$K��/掹A� %](D�R[�\BᶎLߜ�z�?�ј�2�]��j�'g�M.E�����u�FC����|�p2�7��I�ֱ�;^�Ujh��9������H���1+�F;UX�k(�qlދ<�����L;!����:#��WBӠ���<�g��V�Ӷ�壷R%���&�v��`8�AnB4�	��7�_6c��6񨲿�@��qeY��ڙf�a/���������G��&�,��"Dh�ﱎ���m���<@ķ�M�.|��^�A�^�3�4@ �/����E�iZ�S/���7f�]qڑ%Ck�Ϳ�^�����
]u�����o�C;D�]bD��'��To`UPo��bӥ����& ���	��*�`X��M2�5�Q?j{@`KC�9�G]��C�N�r� �lA�R�z3�9&w����@�m�>�ɮ��V��8�+���n�!
��}� �	����J+S-�����l@�b���<��9~�~�1�S����/�2��C~k�$�@.�o�RNA��j�{���k������:�f=�n4'e���Pv�y�PF0�� ���3��"�$6i�*�(I8�����e"�Z��pg�mN|J�$�	y6hp��ot�G�a8�=&@���JI���F�5k���d�$}d�̤ŉїۍ���v��~!��S* `87���������Po,�vCA�s�g1�v������W���P�
�'xMe�V��}���=ņȶ�6 �U&�eH%��6����5��%5l6"�deuO~R�R�ym t؆)�#mv{!�[��XcP�/��fG�����
bϠ��@�k��Z���5	E��3�o"���W��=㇪-�n�u)��7D=	L���@���	�@J��g�<�^Ϫ���s�?�C�SJ��o]���?��~=�
�	�uߦ�����?�@k�!!�,M�z O��S���J���Z-m��ô�J�[M ��\q�`W+�iV�m���~L��"�G"{��m �LrA(�W°��P��
�y5�oȃlz�� ����G� �b�xi 1n^��7r��:LȦ��!�J�	T|��͓��"�����Hغ�o8EW�������.�ٛ��u�z⏊���l�3�D�`��B_�<W1~�Se���������M>6|D�~�D|�a>�1e��#�3G��,�)���W�aW���陫���)�1�;�	Ʉ�$�rJ�>��Z\�w0�؁-0F�f+�P˂s��Us�aY~+�w�/��tBM`bkP&���	깊��0K��2���#U�dVXYHբQ�� PD%������a��K%�2�	^u"P���6��vq��_T^�?iT�������n��gƆj�M6w�e�V�~�`�{�$_i��i�K\�[����J�s<"{�q���F)��Pd�Mg'A��m:'�!�ǡj�g7����s����g~1A��n���A��ZʂE� N?l���dVL��?�ݓFy5��4�ߑ}MY^7؉�N��ܿ #����D��*�96�!����b襶e�(�
��a!*���dů��M
�b¼=��bx(y��@��K���k'H�w��pO�at��;���	�;�L���3���]�j���Ԇ���d\�N� v5ilDX�Y
�!��o�C�s��[9�<GGx�f=�C�]Q$�;G�*;�]ja�s�䥳�1h�}�o�*)gxJ:����<���Wɽ��ѫ)ӎ�$Me�Sͬ���e�Z���B�IB�6.�:�[&���3�$�*�g똙^�o#z���s�k;�jH���R|)�y���65�l�#v,�f��1}�-7 *#�$��8���y{&j�g>���}��sD�{i��X�3�x�M�,��5�w��'�>.%�"⌌��BG��Ovz!�+>�5+J��l�������ć����xĝ����D�/{��?��|^�`E�y�?��`η�+�)�U^����~��G#s�a��{�D&�lI~���.́?������#�m�\�Ll��^U�CB�5��4��6M[��@������!E�[����f��ޙ�+��5$�^{>'3�A�?�.�7�	�8����{��d��E?��!�L�S�/J&����;J0����G�������5����s�۩_�3Đ���D�}�[�H�詡��&��O�>�ϽB���liͺ�_l�-m�����6��/m��'���D_&߇�w%>{J¥S��՚B��i�-�����v��,��ҿ?ߢ��F�v ��L�z`���5��S���򕪟{�:����ic�����,�ߋy��� Ԓ