XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���S�)7��ХBq*��*m�@��#�j(6Q��R���B�Y`в�w�e�ΡK��T�me�@��mW����R�e�S���� ��@�>�姁��r雠�'���������7� �y���pI	N���M�L�.�R�} E!2<����*�.�~f7I���j�2���]��(�d�Lj��3��4���mpQpu�ޔ���[���E����`�}��
�3V�?{]�v���ҁ[h-C������G��wb'��n)d%��"�Y\o��	w��iV ������
�#�Ό�A�$P��:�f����V�M+}�@5���롊�v�+�5k_��M�X�v1vzf
�d5��_�������*=�Z���<��(���4*�T��gPJ�%��Ns�1�j �R��yZ�c��d�qro<Nq�4�����:�g���K���`fH���`�R�L�����^B�4U�p�F�x'�v�)�"��9A�5�-,�g��sӵ�Yh��%pNՌyK�"g��|z���3�r$6Ęw�?1i����yD������?�9�xK�Nm�fS����5O�d0��W/ɛCq��ʶ�f��h�P&�2��L��ɚB,�w����x<|˸j.��2	�럯h<���ݤ��+���ΔlJ�J##�B����q³�����I�Y>��yx4��֗q���
�������W��˘2�n_t���*�3@�.�f�3K_V�\Y\>�g?t��s��3囥�v
�Y����XlxVHYEB    47e6    10b0� ��X���H������s��,u�:�$P��*�^@h��b9��9��-J7P��lz���,_�+�v���2#F!á�?a��Ie�unKT�b>w@�*���\���|�~�<���_Qi�X�ͼz$���+e^W��G���j+�V��&���j#���Y �� K�����h�)��%��f��c��Y���c,:q�$�1��:�k)a��}�X(�b	��8u��˹����{�_�'��F�GR��ȁ���p`�hj�b-��������>?���^�
�`�~�+�_���!$.y���<Ivx���ùhi��N�������Y�����$Qn�9G�aO�W������N�(Tg���v>��G�,�&�n�����/�S˓(sc�����װ���~�B��e��4?$Z��A�Xގ�嵚�V28L��2|<�����k�5����5�^AgK��$[����`p��'[�oY��M@ohe���-�msnCwg���.8�/�d:���nN\� L���i�ݱF<|{ņ�x���F���7���o�%����Ma�Rs��@��:k���������<�	F�{�*b�dp�Mw�c�e ����y�I7$S� ��ˠ�p�-�����Y��E�Dމ�`ʕ��T��\�O��,�HP��N<�����~$.L�?/���[�I�o>H�&���D�|�G�1��l��=!Rk�**f*k�N~q��ʡh �(4m�&��P�2��B�����Ԩ>r�PR��2o߱�/�f��!���hz�{�=5݂�lL�X��d���u/�.R6��T����;<�������^��rZ�[ƇX:�9X$�ʯ��0:ʹ�F����[2���Y�=~�����8��:]hk���jB�R�א���Ng���j�����Rd�gו�+0ͭЀ�ܳES�������h�{&�G"Ց�U�Z2�y�6=!������I"G������,)�N�Ь���K<Bf��VN�$�]7�A�<�K+�/I"����賳�,$��ͽUþ]<���T4�/�w#?!���E�oTYƫ|�L���u�����&Ig������y3�~��r'�	ʑ�.�I
A��
�=RV7��5j���h��3
@A�@ �՝M��7,�YH�)T`T�6ZK��kx
��x���ѕ-��#0��JSӿqH�[
S)3�i��'�rh�2WW�\�y��K !~�5JN2h6,
�!�����˦��2\��0-( i|UԪ�(��	�,�N�/�ѝ{�nϱ�U"Kd�H�+TT�vm{Շ��Zp���v�%k��!)�wY����o	��*���!F�4�ɡ�D��7������!��W��cm�zhq6Kv��@���1��h=��K\��hZ#��HV��f.���(11�1��s�B!?ǬU�a���W��UF��/���[�LW��)�1x�f	�i����/���`�C�aۭM��`|�����V^
�2�y����j b�PF���ؐK>h{�g��k��.�obFo{�;U�F��݊��m��EL[�5ҕb�É����v�^Ɂ����Z�[KDP��5T�:��>��%��:\�3���;�s�#9�7�pp����# N��iԇ����~�)�c�Z�Eo[T���d��j�U���b�|x��=�� ��:��%1<�Z����	a��(���؏r�'�=�����S���V��J,��*��6�4?f�o�I�+[�c[�Mˁu=h���Г�4Pھ=tn� -=r�{��brpញP���7W_��=���6�Rɫ���X���v"BO/.5G��&��;�w:���K*�Fҁ�V�lG���6S�3���SR�S�Lbri ��5Nb�{b Y�B�o���6}�f-Ю�_&N����r�w����VF���'�k�[�:�
*�2�֙���w�E��'2��Z�P��
���|W<�FN�{b#����ka�zL��Q3���`1�# �C`�G������w�,Q#�eƨ蜑�]��u���)x.ƪO���i���-�Ds%I��;�5��2Q�$A��U��%<D1�����d�B�a��fgŏ4r)��!o�2��k���G�A�u�*�/�*z}?b.	Bg�o.�ǰ����d�cP���Lq0*��b��6��O,��D�������K±W�E'PFƨ3���43��ԇ�ʯJ�IĜ5�v��ı�9�P^�$@�/\��(ƌ'�^���Xt��ȧ,5 �x�ѓB��!ugiS�n��`���|�"�3{�fO6Dv�I����Kg��ɰ2mll!�Y��f֜#��x�mU��e�&�&L�a������n�/^o'�LO�\���?�������i(��t6'����.bR�b	I�����̲(��~��m�/#�B��<���ϋ�����sD��s#�0��1��F,�ƺ���cVJto<æ��Ǩ3�*u�,�B���u*�$f�m�����*Xu�	g+��D��e��]�ˍ��z����ht7�q:L�U�%��͏�r%�{;uUL���T^��#-$~u�]���j��	��'f��~�$ߩ/�\��
/#wU!��55�� }��<QSqf@N4N�{����a8���l�m&�2�A�	���E������g��H�L�L���U#~ʯR�i��=�4h��ħ��/vju�(�a�'�/���,��KZ���A wݦ�r����Ǚ�n��Qہ�&�6A���l�J�m�j�g�f�th�f���E�˥9���.�����(|���Z+x<��w�='��3[�9�=�v�Ӹx<ڒ��Ƭ��ݔ�5��j�r%/3<fK��%QW�4S`��C���V^�`Ts<%�l敕��y��ҝ�!�AS��ۈKE��u�M��7�NsI|ui?8��z����?�S����a��i�4��>/���i��E��3B����m�-�X���8ǰ?�n���u�d�;�hwP��F*B�p^R��9�Ƴ�	��;���G��!j����V��)G??�t�VQ�'��u��Փ1�UÔ	Đ֮c>�ŲG�Ę�Im&n��'"�%1�,�J�DiT�ϑߏ�e[��e6&�#?���-�6��n�a#��8��Z3��%��%�p���b,�����Tj̮��vU��ᾎ�{�f�qH��2�G�3AL��n��n�]�.�kN�E�˒����{��ҭ'�K5�7��R��:T�:u�J�����q��vQ�����Qʠ��NLO��݌��؃�B���gy:"�H�ޘ�Ԭ��=2�BrN���O��nb&���S���i���{{33�n'?屟B�{��y�kn�a\Ҳ���Cu��Y[��� Խ`'��5�W~@Q�.[�s���}��V�쀶�{>��5����.�ry3 0Z
�Yb٨T0��sjs�%LݵyH��F�?��Q���N7W�`Z���pzH��ˌ�A����*�[Rp�2m�D��n���kN��)=�z���G:E����$`XQ�jf//�{� �� �᫪�?�5��*�����(��V��J��^�li*��S������1�(��"&b�jJʳc����	E��U�k�C(�><cT�(XRז���`)�
u�S�_ƽ������6/X02��G6��5�k#��+~�g��l��t74l+�\���΁32V��u�qzf��b ���x>�"	����
nG�أ���T�������?WA��)EP�$�+AR�s����t��J��$\�#�!��YX�����f
.���=�Q~W��!�la(�0�d�{�����r��Vj��� ���1��9�$�[�;�B��X+�(l�x�;��z���e�ºQ���O*��q�����%� �d,�J�m��Sb1�F�r�K,j�f�[�ۂ�K�R���je Y��P���PQv�^ӭ��2E��#0j���^%�oR�{i�d'��S��p�i�@
��Xe�6�h�U�P{2)
�A��1	�E姟Q�,8��J+I#�{~?��P&
� ��m���R�],�+�"�2o��$�D�a���	A�I��*]\����	v�$�*�Gn8)��ȭ��ZL���[��v��%�b�*�2o���I��ƫ��S
G�0�lcr��<%���nXI��T+�Dc��-˛�