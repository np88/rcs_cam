XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����?>���wy2���Y1�+d�&0}Q_n���_Ε٢��;W�.��mM0>'�����ɢ�qZi�9Y��	�H:�6p�Q�]!���_E�G��H;4�(�ǎ'��񨿃`<%S�_u�H
��G5�(r���?��_Dܦ�F��%�nFz0��Pk1�;������Rw��sU�s���OU#~�0�u�7
¦����S�qF�Os< �%z��6��,�{����*�ҽ%�B����:����r��Q\��g�2o(?�����
�QT�J���p��GgQ%ƛc��cWJ����癘�4�ׂ���K��2�qTكbk�vF�04��^~p^ B%�qݘwܡV^naS���<$����\"�v��������� ���5���A��L�J�x��:��X����T|d�pU�4��P@l`��)�p~v{� �
/��bT�+8R�[�d|���8�H�La�Յܮ5�xy��T�K�a�Q�k�}�Oig~z��I��1�π�H�0H�iC�[�A�{� �6����VzwR��4! ���*�n��Mg��l��D��![�+��|�:r�ߜo\��T�i?�������Ƅ]B��4f�Hc"�;�{�En�wݫ�5v���ß����	�ה������Ыr.���Fy"U,�(?3�����A`B����h�o�7$����^<�|��D= ��o�����j`WEpzz���j@o)^�ݯ���-FB�;��O��^��ײ���
��,-�[
��9��XlxVHYEB    8e9e    1d40�vg�Oڦ�`k��Z���$����4;8��)�1Oi�I�R�L�JWݍq���\LT|U|L������Q���� G� i��:ᶝ�ia���t���!�!X��	�|O�mA���5�����	�2���)���a{�&�to��ɿ�����[`Lk��d�&�T���Z�{��1\R���Z ����ăb0)O��I�I�v
pe��9���Q1w)`1}x{�;S�Z�(W�H�SG8˚fk��q�r8v�r���k��J���yF9qdK�[S��`'繿bj7��wS�����W.S5�i#X��?��6�Q�p��/�����;�}�%h���\ ���Q�3�*�kᳶ�Ϻl����i�7]"C����ݓ-7�I���`u@r@��{���%m��Ԏ4Pg��|����b�
˨?�����FD9i2��T�{�񗥗��c��CB}�-��@�`v����F�v����ae�/9�K��tLJ@�} T�&���|�`z}]#�гT�V�B+�"e��:Е�g\{����YKh�Z��l'rЄkqZMeՈ

���c
�7��r�
�.�
Q+鱖�28�5~~?�� ƚY�G�F����2D ��H�]�5q:�|XK���c��y�{��Z�	����i~O�C��0S|;�����7����[�d�"m�����#}kl�A��?��
b�Aߣf		�GUP)��BC�c�|г�E�ᑿ��D����
H_M���	i�\�p��8�0؁?<�]w����t�7���X�R֞�si!��:^����P���U������}RR��^�[�۰3���yC�Jd7ُ��3f�_�Z��m���q�Y_��h��9|&wv�DS�87����:^Zqy�S�a�q���ND�
x�,[��YT(�^V������;fr����*Vנ��Nޮ�@u�|2���\�껱$Ʊ�
O2e��An�V�]��M��	m����풽Ĝ��v_f�\%\�k�5�;�Z	��=杣����%�9��@%y�O���z�N��SO�a���<7��1��,�}<�ԉ��E�idc����%$*7{oӎIJ㓼�=Z$���m�{# �juL��H���j�g"�f�f��^����8���˂gl6Q�B�%?\6�Ī;%�y�r'@��>Д�%Q�.H ��;&�����u��F��AF��� f��?on�-I8��o������5��8�J���3�ڥg���ϫQQ-�v9� ��^�RǏ'�a�*���q\S�iq�W�`8T�'4��M���3�up�X٬T�5�����|��RП�l�
e������f�$$��䉯6���L�f�zy�eВ�oF��f(��b�4�Q�}'v�=��SL��O�.�#���1� C��JN���Y��`�p�U��z���������&���*�������_7v���=��B�
��ݕ��ܲ�G��*��>%QI֕إs���Ĝ����}�:Sݔ�b��V^-�8��9�W�*O��؆��$ϯ�=�s����g�h#��{s��^_��ڋ��\~�x,4�"��ՖS��1ǯJk����E?�\���j5�6�E̿-��.�lH>���G9Q+�P�X�����T B8E���LUB��U�&MD-�����βY�4&�Ä�a"����8(�V�������#�g%�����ǇQ�	2P��)M-r�� /r��vC��O���I�͎�/	��~�� [��dV7��e�s�d4�`\�����>�􂈝P���H�?*쑨��98��}�ћ]t�ٙةU�Z躈�K��ւg"�{�O�����;�t����+�|	z�hr��C�-����:]�·��o���Pq5g�(j_�o�a?��g��ںm'�L�l�q�QzG��o�ۘ�˅2>��"n��Q|�0�m띴�
�N?;�D*�pjk	v��8m�^��9|�$"ڕF���:^ ���&�w�T��a��Ԉ��(
?���6a[-$�
�[�7r�e�{����=����X$���@�q���A�`g���4\�cj���j[�,!{�
.UH'�[vB���o��p��LXé��[ B���DC�-�f�j���(�]Zz����NL�|
������Ө�3U��	XmT0�ta�hK�ܤ�r�i;�M&	6�J�(z�ΔS��-�6�)���ҭ	�j^�Э־G*��9z$�ޒy;��{��K����a �3n �*YXQ�GƓ0V5�i���yHa�� �X�^�d)H�5�,`Z)oC��E0��^�V�M��sC^S�]�o��κ_�W�^ű!qz�7أy3(�t�c0Aj��>Z��2.�}�aU�h(}��]!�h9dM!�a�~<\/����_���xjz,	�0���p3�U:�,�~�Ch�����IF<�5�L��{�Z�Mo`�h�6����58�s�1N�}��]��\��wп���Y�]?�<�/���+�}.�b��OQ���yY��M!)�軇~*D�S4����\|i�}�**|�!*�P�B��Q�q�����v��0����[➭̧�K�!p4���1aH���=?h�@{�:�gL��3WP] 
�H�8��3$b�m�P$JY�Fh��E�jYӻ!���w*p2�`҃N��;�[�I,:�[���P�"�d����(��|�#$��LN�_��i��o��K�l<I��T�z�ژkd��\7���� ���2����8��cjN'"}}z�^���d�6H"x�Ln'���j<�
YD�B��خC�ߡ�����0���̓m"!P��B.���-�T����LGt�?ۅ�.�����۔x����(�a"��s:���nķ5il�SV1���N�-�h��xib?9��7X	�x�Ki������?���LR���k)�5�;Y�X72Nd;3XE.�Y�w	͏Md�1�fޑe�I��,�E+aM�ު$�N�bSn݌F$p�"��������2����]7�Z8�H���{�N�����1�+j:�=N��.��E�
����g�Xl|��Al�8���V�K�[f��jHCm�8����b��E���s ������� Pe[��2o��nűnRk~��U�-�S2;՝��l�7��]ӣ�D{3���ء�������3,�@]�]"�PGю	���^|�`-�� �ڊZ�Q/�7#~M��KZ4�g�j�������\	��	v믑^��onȿ�g ��u��"�N�[S՘(v�2-��s�BQ܃n�M��W�i� ����-���ں�|܋>Z��H~߅�4&��|E�q��Q�[���29�x�Z�X(���>٪�xc�vnY)�����㑶���2�Oox
��{fM!���H�,�;ӌ�ց�j["����\kq���-,L0Òbh\bhʘ����#����i����B��f)(8���}�O����Ý��Hm=�08/�n��i7޽���] ���l(s�j�Q��R��Oޥa�c'��S	�������f� �[9��YW�Q�� `�%��˫VT����T��(��|i?�,8˯�^{�g�2���m��s�#����ݷg�l
��� �d���
fϔ�,���Y�X���Y��З!M&�ys�U%�(������!��V��4XTF�N
@ɠ��d �[�]�]�OH~��z`I�?��8Kۣ��|�x�����A����G˾�B9"�=������X�P�u��d�Y��b��g���-�\|��t�J�_͙%
T������^؁�?�#�9Q��dθ���*$�"�Ϲ�0u	)���V�Lt/z���=S,[ϕ��A�c�_n�$&��3ZX�1�(94(3��k��rv������{v��ij{Bm��.*�j�F�F���g�[9��z�Z	s�Ė��BQ?��v�7���.�[�*Ӆ�ȯA�[��gƟ�Jn�����K��j,{�lZ��D �w�504���@ͩ"�_�6���}�>�-���'���鯍?p���G�*z�:b��`F�������^7*2ǲ_M���ǥfC���	:,s�E��	�2���V	)_�ތ�i�I X ��| �8�TQ����88������h�F��O�Q,��F���]0l)�R���q<��1�.Z�L�'p�,��T�t ,�xa���hw^+��g���+���=����������.;�?y�ꍏ`���;�˖g���'%��6eg_9��D��c�� �L����V�ldڊlӏ���&/�� �f���@V��s^Nb�oi *�D53��"��;X5E�`D�ީ�˦�>���"_���OZ�8�ŜOQ��R|77(}���.�Cx�/���4h9l��Z�Ipfh6�A��tP�CxL�C�4ۈ*:�\�Ο}t�pv�M��I���^
q��k}�n�Z�;O'�φܷPt����O���sQ�з�����q��o%O��DA��ǖr�k{Aw���U�Wh:_�QI0Zr���w����Y!������G�~ Tժ���
�����NֵU�@+J���h�X �H���qu�)�~pG���V�l�ٔf)��1�e��T��sW���%�h���ŋ��!}�z�bQ�~�n�XXy���b���B�9������d�'䱟�#�m(��}�<��&����S&3T-/x��`�I* "z`:w�U3$�%;R��]��,6 �W��.�E�����&'��_�#�MN#��~a
�q��f�!�'�d}r~F��́�<����`��L��״4pKR�&BQӠ�v��!Qڊ���WD�o�N�p���������Zd�@Ugb�0�B��܉�E��ڔ��j�HN�>�=�&6m�ܢ6����ʺɌ� :^#Mmm�,��t���~��_�ɺi*g1ҋp��ҧ�x}����p���i�8�8 .7�Pƈ�-��m��!t���Cq�	UB��)�7����:vǟ4�Ir����9 �2F��d�UV�2x��o٣�/�ڦ���ƥ�k�:��~y`Y_�k��X/�'o:
��BtiR(w*#p�������oa�Ih��-�F�b�*��B�'R�{qߋ�Aq��{+�JC�/(0��5U�FOG��	惘i借){�A�]Ϙ\�e�UD]�Rܱ�djz�p���*�,Lu.�J��ͣY.Aτ�f�����X2��j���t]J�{�&��[v�P�=0Ԥ1��,�@��(���8��wm"w�wn*N�����<E��l�D�+
��Jx�
"�r�^�J�#O?�d7�@3*��.s��7KE���m���E��g�e�3d��%0�n�B��q4]�У�y]����w��GNӊh���P���y��Ը������}@%�\��ZZrp���<5�V�o�ZG�	��;�i=��b�E�ly-I�m�]O��BE����K�hbR�>��oR�%�������]��y[m�d���ȭ����(̭�{·� Z�����֜�����(_��%�ġ�*� y=�b�:�z�.]�vn��9������҃�6ېc��jd�"�X���<�T���ݺ��"N�|h�ZFiPWɯi�I��e,�΅wglm����NMI?��K�u��/{QJ��q{�Ρ=���#¦A!Eԗ���D<o�)Q�jW�x�^�����"?+��}�#�7םzL��ZsF0l�����̲��\~��n���L���(����4��9��E�Oc�#��^yD��{�%F�<�)�!0"KU~��
��:c�s�4��P���Wo!�>4Z� $!#gN ���-P�ĴS/��� �斉n����2�ew�*�o��ؙ#��Xh�wդ;\!3�
�yF35��)yn41��ϣ�+᩻���%�?�O��eu ��ѝ iS�ʉ
�{p�^�\=\E<|�%Km��Mй�ѧ]��W7rjj�o=�֧?Y��{�=�?��H]/h�`Ë 7F�F�9Z�uy��r,N�y�娴a�Y��g	I�}g�%S���9l%�K�S��ƽ�� ���a�$���2��.j �Y�u����n��ι����O�3GB�u=V�SbW�+?0DH.b��f#{G�k�aN��G�p���ʁ�k�uY�;7��8$��m ���Ԏ{�X"�gs\�M8o!(��Tl���4iE�C
 0���@���.P�L@tdq�.$!0�#�����t�b�oeU�Z��i@B�.|y���rus�NA5-��s�d��G���vZ5�)�3'��I���1E���v�	2他<�nMŅ;~r��&"Ca���[��9��BF� ��������5���!���Q�,�rt�������\ܥ���.�	:��#�&��wHG�nsߢ��yq��@�P��Y����G;���4LtuY�ӡ�Rn]��4���~ g�q��rZz��h5��wVً]F��4@a��er}X"�p�2�e���J.H��4�Թ9���b�=]נ������{Z�&��<��?�+P��p~�3�B�, �ezJ�7�[�����J
����Ľ��Ek���+qE�+�#�|4�j��4BaUOg �Й9'Ց��5h��@� s����BÞą��oJ��%2�ʨ#)]x���2���m����w�	����Q6[��X�dh-]��tj�B�؈�E^���*,r��m��(y�XC�H�(��]���3Pɗ��RPEKA3���qe�u����$�;c�p��Y�c�"WM�W��v%1T�}W-��j�O+-?ݔt�Ʀ�DLm�r~��ˊ��5��F�Wk�H7saL����Ƶ�=J��ٖ,5[5Յ�q�ON.	�0��
|EY3C҈}��)�3_���2VR��F������d�W0~:f�n��-�c�����:#c�c�y�h���T����9��4��m�<��;x&�i��nJt.�A��W.i�ʅ�2�m!y��^�����հ�jZB�ɞ���n�}��2�g��ʬ��R�Qa��3����))T�/
�1ՓT�>tZ��w*+~��n^7H��J���/^��˹	���|���y.Q��Sɋ��ոPFߎ�����{>�%0v󏚞�@Fx�u�dƧ���+D�݅G(� 6�6�?�'�)U}{�kK~�a&u��e!°�oY�3�(:�"�.n�P-���O��7����?w-R]y�o$J�2`l�	��"���,_��@�3�����E�p�s�7�������1)T��`�Ղ&KF��"='�V������g�!�CV�c�L���y��P.��k����|��*z��ɼ1'������'s(��G�,l(���"$�m�A��On��^��"�<��+{9�d��V�U5������}V��<��vUjءcwV����
