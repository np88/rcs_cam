XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����;��Ёr�=m�%���=�1��M�]l�*2���t^%
{E���b�����hh�-�(��VI�DI�klMx���P����.�(RD�<�	3*�҂�<f����B�-%�`;#�"iP�kW+�+��Gy�.��g�v��9��k�+ Lx�#�j��g�]A5����G ����SA�{��_��Ƹ�6@[h��Hq�?@�L0�z�}�h9�蒆��qJ'��0z�2zې�%�>��iMf�Nn��<��/�@�4��v��ZR�������v-�Ta>l)(̕dڲ�O���2&bU�%S5o�ǆ�'K�v������C�����o�/(F�B�֬�)l�k��Q���p'�+P���*^]��VgE����r��x�#(��N��UE}8]qڊ!�0�^!��tjY�˂6���<4��i��?F�S��&}t'�\nJ��t9�����Nxt��|b��Cx2tG&<�'�e�^��'M�Wk�0	T��F�a=�g��H��G��$�I�d�4��"���~�T�i�}9���Ŗ��\��]��1��/���v��C�jx�D9jPD�(1���i֫%դ�9̙�u)�	K���R��� �t!r{�� ���+���Gq3h� �[��Ǣ���s�T��:�L�B CB�[�/}rA���S��&[l�uew'ۅ���3�#�(��2̯v���ɨ�(��*����*�ݦV`��}�nHy�:Z�w-v�c�\�(Byޠ�c�r�XlxVHYEB    29da     af0�0���	���.{�4sA��m�Y�8��n�a�MQ�b��VɄ��ذ��T>���TUS�RJ���ʬ���"Z[�+4~��@�Z^U��T�|��*�������C<paR`���������y��<�_�����:Z���u�H�k
�J2<3W��(D�Y�|��x\��kn�oyށ���߇�[(����p�4�N|G����@��ȿ���}��Yv[DE���̏_�G_����3�� �s�B��Y�J�l.�_��!�u�yx��	R�V%b$ns�d��=֭������/5�G����5FlG�oj��� �K�Z�7�'���䶤���i�2�m��=�'ۉLd�e]_T|���h�G ��Q�꫘~Y?Ko���S��:���h�\R;V�ei4��t��F��N2�`ԫ^�ۑ��0�6�S�(-�T<�
H�W&�=��eK0�S���5v�@��Yd�g
����Ҟ��-u?�U)��uvz�6�j*Vh�YAl�qqW?��F:�,�"!ǟ4��$>R쯇M���@�~�$ҐWv��X���� �� _3Y�Ǖl��$��������������\�7`���:�Q�Ie7�5D|���տ�冒u-��s^f��L]y��G0�>�VR�K@Jph=G7�B��k8$�<�>K������7�B�f��6��T"�a`��m�@�����M<�r�����̶�R���
.��*���$�\ζ��aLs$�B�>���nt\���Sp��,4�yY�������\R�}���{3C�J��L���$�iT�kҵ�Q��O0+��<
�J���z� �R+c�=G�U�Yt�QP���:פ0s��=53Z!�: 6'�G5b�C��]2-�7\�l��9�&��^:% +,����M�ދq��b�.qS�pc��`�� ���*��,}��n�n����J�׆_%�����KOG �T�� ��3B-T����]���8����䄐��7E�H3���D`����bK=�Xf�u2�m�"�ǐ��]2�j�&�iP����zz��ٽ���T�X3��ӝ2ˌ�{�1���l���W�%u��#Zu����[h���gHؙ��N���lE"�E����^�6�B|��KQRn���$�BC���a���ʩ ���*��A�37�@<z��O�/6�}o�����4>��V������I�a�\,��yA̎�)��2�������nPj ��\��egv�5>D�K�bɄf5(�i�O��Bs���A3j�6�V��%�H�I�H:*�;�DR��K4*zs}�4\u�����H�6%����� 1h ���|��(gq��M��֊�f�Hib֑VID5hA{7i��J����C�WB��/G��B'�.�m,*�|�!��l�������谴.%�Z;5��X]�iXPX���b��(��
�k���4@�ע�l�im�M<�d����3�nT���JwK��o�u9�"��c+�1 <l�m���R"qM�V���ߴKR�Z���/ߏW���?M���,���r��-܉�6.w1F���H(��l���F��c����i+��қ7$���I�C�'��1����3��S�;�m9�@��d���є��n�N$EU+W�j��OW7׺䑔�؟1��T�g�"'�� �/";R����+��eP��X;u򮭡���5ZpmU=A�_�U�nt]��e�y��0=�
���/ݸёDf���<�r�u�8m�ͥ#�nK�����2B�K(�y� Ə}����5q�ϐ]k	/�+#���x��^�����-���D���l�V�����E�����/���� ]��E��4y�����H��\NBD�F���j@R}�c쥺��l����_]h�0��R[�QO(L��%&�'�7+�3W�"l5
��_�uN��1�CV��j^?Bn�c�]�*y�C͡�!�K�"AQ�ؽ����e���X�
�3�OE��N���Yۘ��	hmK�	�H{{��\��>�vD�F����o#����7��A�9�æ`����$��E���!L�-	T�E��H, �\*�=j"r};W.u5�����c�u(��E�B���X����t����~�)�W��GE��Н�"QW��B����=�`�wg?Of�ⰶ[b�Zu�>����7�= �
X��q�>����d�K��D�Q�B!�$&,��n]@Q������q.�t2l�S����]���5+�3U���\���'�4M�#�k���Z1�n.�8J%�S���)��i�\ q�4�	u�_f�*X)�f�p.�A�k���Ǻ�{~�@��HCY�ž�3D� L��Z>��dު��<f�U���l7��X�cy^-�-cW`v�pH���ŀ�}�#y�2，�ɂ�aH�i�����[R�/M�2U���-�ҵv�w��͏2��L9�{��MIFQF���J��v�ÑT�����,_*������P���c����	3{�mB��nqb�M7�LĊu̚�֬:u�S�����l��F�:�BT�{�>����2��&�f@���F�"#M�{=�w��b}'O�``T����B�}Z�1�ٗz=2�#)J����������;\�;��9o)zz�;,7lU��:���wk#��L1��6�ӛ�ʊC�ؾ��$w�f0�`�c������da����=P8�������x3VE)�y�EsS��@#�+�H�|��-��JFUn�&��g�,\[R&_R%�(