XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��$�tkJ;�N����B�5�mR��ċ���}�^�xB	P�n�YO�����xs���3�$��PX؈c�8r��׵*��W�841��p�b����]�Ye�mx��	yd�J��L���/Si ۧ��c�j�^�_-LD�̻������ �PR)v:�sm�&����X�k.Ͻ��A�ܗ��G$j4D�L�9���-^�8�AW����e�7�J�	.�
O{·3`yQ�&��msy:G}A����)ME0<������bGO�A�^X���!��	-�	���|������Yp�>oδ�}��|�r��-�|C
�ψ­&G�$F������$���A;��bz�Pl�k�\a����A�0���A�����%����:���:�΀ݮ.���J�
l�~��L\���d?�e%�����������}u��$��d��v�+ï��!8��'Nr���{j�g|�P��g�4F:�a4Q�mRa��d�]r[�CjF��[�%�Q��R�.5\{�z�'a(~!)^��ʮ6b:�e�Yk2-��8�5�; 筃�����sp]&�e�da�+�9]	gY���<~� 5�ϲ���� �g�-9K�R��W�Y�8|קG=Wܺy�u_�f�|#���Q���_�̧Fif���x�g���E_kH4�QA�hl!)�@ }0�� ��f�N��(�v�l�5�5;JJ�A�s����vY�4!c�W��":еБY��['
caY�>0vYXlxVHYEB    fa00    2900�_��djjnq5���Ԕ��i�)L�������1��������ՓM�d�+uq{ٲ�#�[���T>���[x���WgH�=A�Sz��v��vqݍ$n�"�W�N�p�ZA=��j!�%%~���������ի�`�r��Ϋ�LC�n�����%^4(ƩR�O6ȓ����7U��/Px���ɢxB�R����^�n}l��;��m��ic�v�o$����z���4�)��ގS�
u�( ��D�"HS���ǁ|�e����d�U��R�J �g�'Q�yI���,b��� �?O!K��'�hzw���;h+
r� ��g ��:F9��u���l�`��f��"��>\�	V\IU��2�a�4M��ǟȉ��@�r���L�����A�W��0�d��������>o/��=(M�w�nE@{X�ʧ��0���ގJT�V��hYI�-ȳ�m�ܽ���54�s��v��[1���5��fҐ�a���%l��#q�����m��������00�j����9�@����#l1]a���M� ��1\���=R��#��C\�Lg�lz	G�'��.l��wvBl�;�>�M+�f�(��t�u�*����T$�	���y��sl��Y����=��:\t��Vj��N�ߵޖ@�M����s��in=��������dT�+_�bp�	�	�S-�g�r��6���C�#�M�}��o��� �~� r��W�-����p�e<*K8b�&mr*�W3���)��t�^EQ����pf!��|tc���,����v�J�S���\@l��-���౵6]Ռ�31�T$!�z�b�!�`��1�?�8����>���Ֆ����2�ED.��ȝ��=j�
�I���[<�=�'�����6ۂ�����A]��ՁsH!x��<�2���.>���cА>ws�U��Ee�Z$��3�3�K�M��:�c�I�Jq`ϞRo�A��$�)�c\ӱ_yV�%w�v�t��j���!Tl�dB��)��/����R}�!0b��(�Ls	P�������;$Fx��#��p}݅�~Ѫj�;n�%[��M\+��ߛ��ǳݣ���ed��J���Ї�����7%�(z,���e���x2���J�����uQ�-:(���è����%��bxI:�F7�ڴ��s�c�8�HB�]�1�����PӪ��H�<;�$�O�&��$2�;
:��*U�Zh�--�M���{�ތZ��(T0v��Rޝ�ia&/��c�}�cmA��7�I����
wj�BX����/!�e�.Uc1����<�1�0r�,��c��:N����YL��v���]:7;��?(^��?c���Tӳo/vbwe^@k�f��6�#8��@0�4JH�^�&�gT�������o����Ԉ�,^�"N��0�"��p
�7��-��	�@9�t�O��ŝd�#����So��>Ym�Ɩ毇7G��>���H����1���*��C8��)O��~� 0y�A�A������t��8X�D� ��4�&k��XuM�ߥ�5��4Ӄj��,�b�lV%�}�gt��c*α�а������6��8�`pg�1�x�=UErL#{�������%|5�͊OO*�G��>����.�H7��HΛ�/�"&u8��Uq,�Y��)�1fT���_��Gj���l5�r������lR�Xp'���`����� �\� 4�W֛	%;�\k{�F=�Y �"s�Nnz��]��C7=�0����5����9'\���Anlw�w�T�LaG����җ�č�11���q��  Xh&n�`p� Ǽ�Kݾt�[�`O̒w�E�J��#��@�%��C3�V@v4���d�|�(4�*@��6��f�����ʂJ2;x9�=gPյ6W���%�-�,�e%
j�휴7�'�ۡ��,My�NSB&V�w��
T����٫��v왏2e�"��!O��T����wf6����/j*jҮ/;�$|�ES��^x�13{	�?0��K��S'�c��}$� j!�N|(rֳ�KQ�V�\ �O��F����J˿N��E�&�AXd����f�Q�J决���ٽ����%��4ţX���,1���n�ذoŒ�������d������q�����9Q�}�)�A�8a��Q�4i��d��P�0u-�Kn[�Dz�kv�F-�kbz�eH�c�X	}.1�CV�"�3����)�ڃǷ:�d��=oQ�Qcp�0�j��4�{�7�=��f�3���:zMě������2�~� x��܈w���'9���|!�sl��Q����k;3�#�T��X�[ʐ 
xH��CJ��{N
u#m�f"9���uR������T�u���kƥ�r�5���4.C���ꋘ��4	�V��L-1r�f&��^�,Ԋ�F)ԏ;����b�O�07s�>����u�Y�����������`N�,y|�;��Tω��o:�6�u���I�[ă?�Ɉ�O�4SA>|h�5��BX�NPy�*�6ғ֢0tC��索(�����w�T�K���8m�n ���ĭ�o��m�W�xGf;� Y-���b���S�f��a��w�����R�{�,��Lߗ�������o�U�)�hxO�O�]g��V*l�i��#���$�t�6�{�,��������
��>="'2�ɝ<l�Z?1��	�x0 q��w�f���﫢 ���}(r)�/����0��-��l��/#��P��p��
��y��R�{�8�!Z�o��8U������Y�0�4��k�9[���ѻ�VXk����)��t���)�Bej��O�� ��Z��؝�'��UQ
���Z�D#�e��,��~2�Y�&jG�sG;�g���e�Y=;�:�y��6�^���2�RF��io'O���Dp�0|��M� �i����G����r&�Z���q	�����4Ue��J3�+&�/�d�EBV���R�|N��ߍ�����d^��t�I
'y��8eU��*وzp����g-'�Q� ������M�����dZ�"��Z��s���]=�y�\�#�g�)I7�ۥ���K��\|^�T������Z��U7��5��o+���x�a镅��Ջ��pܕ�$�)�g��Q&��oJ�?� ����W�r��Z�P�S �B�D�d�МO�r$�y,: �'+R�k�!���
m�9���{ruN��";Cw�Q�邈���@u5$�����jJ;��@BTe�Ij��/��!��Cخ�{ha�c����㦁|A)�C�Yҋ�V2�2y͝b���@A�WBƗ�M��Bn�~ӊ�!>�i����'�p�-��j��#��a�V��������&e�=��`�ju�R� ��jr^"�x-��X,�:3�p�5�dz��|�87c0q�>k#j� �(=�´�ߊa*�D����_qG�%�;)eR �G%�M�g����/�yl��a_%>���������5~n?�-t�Rj��8��錛c�_�Ңvھ����N~�6C� �N�q8Ĕ�B����s�#?R�Q�5���=��.#N"wD�uL�N@�e���or����ͺ�����^G��PO�;��"�\��A�b �r|�O�)��P��%��#t��c�>Vh�;"Ij����K��F�&(F���������;���n8Ş�.���F��U�\C7Y[��6���d�[�<8:��K7��֬�]xD�+�b`o�������bD�{g.�I9)nGe̦ 	_�D����H�H��K�9����R���7i
R�M��8�r6Á�/^�p��q^Fh�����a�{�6�	R:�c�轖RWV.�;�s�v�Ԋ��`Ɠ���	C?��P*'�2�<�qz�VJ���B�t�A)�U��<�7L�"#����������"-�5&E҄����v ^�
0�~���:�$��H�it��Ls7�Y�Яv��;�K��6�_{MA�/+=�Ra-�T^]���cf��Ɂ���9�U(������@�� 'ˈn��E����3�ԜN�Q�����7'�ٛ���cL �CMOl�U)��������fT-p����� ��V�$�8)e���r��jgE�(�w�>L��h�1��H�*K�(F!�?�����3	��7�I�pgXaY�9�qr��I��'v��!O0^9EV��v�\B��̕�m�D�FJ����e�I�L���(��E�ٯ�gIRcķ�V}98.����Z�7��wS�����/�f~��c���(���0��b'���P���׽���}�i��8�Ը֙�1Mre����׀-P�23dL^w	ݺ)<����z�y���~7���[���ji���U>
r�oh�8���+��G6j����S� �DO^��[W��ȥKоE.#�2p��=�(�vU�1VL�����*�q��%�5Zs�}�"��M>�JmE}
�Xj�Qj²��
"����N7�l�d�9o�X���4�CM��]�u"K��4��P�F^�3��vU�?ϐ��S��]gj	�K�T�@w �,|�p�(b�!{�H֪�L�h������k���!���KT�alV-��q�k�b�E/���g0O��[\��G
8��H�qy����wa�By�I����2B��	�̡k���a]#^�	JҖYPs[�K7�0�4R�0sz=qn\��^��X���s〘C�ʢ��U~|";�u^ݗ��I]������_,�.�{��;&�!��@�胫�1���5�̎?��AG�)Y��)lv|����[� �{q�!�1�^�\����Sxz��c�Z迢�葮࿦]��1����sT�g��< ����i�u���ȩ6sǕ�W�ݶ�(� ҁ�£t5��������=�C)i�%Β�������]�G�Q��}����c�ܯ���z�,�Q�OX�Ōu�'����᏿$9r�e3�����t&aU�Age:}xչ��E�_�1Ѧ���['�V�ڔO��C͗ �J��w��U�P*dq�I۪��ՉmQ�[�WBnD�)��|Kg�[pk��ٚFwE9_��i�T��y����3?�Rf[a��-C,��.4���A���q��/O��Z�7n��,K\�4���6��KP�7�&*���@�)��Mh��uH��)�<��}��C1j�uՋ�n�
�_?�f�o|4�n`;�P��4�d���Tг��8��Ja:�D�����c�]$�䛔�>[>!�3Z��!�x���}α,������Y��L|a��>�o$?�ZT��^�B�x��Ȁ�Y,�R��	�	��Sk�s�x�0��$���Hpz�ZK˪O`��v�O�Mӫ>�S�Ɛ�s��Z�$��zD��n�����E�ɛ���x���h��oS=��⩞�o�˔<�i��91EW���F���c:^�+#sQ���$Ϙv�f\��_�Ip�d�Cv�&vfd�����J� ��L�>#����~2�����)�ƛ]z��,���k���}�F,Cm�g���΀ް�IAt��eX�H	L���vAN16q��k�6����*s`)��#˳4���A����YŕR��c\-r� ��dMjL�����2K�/��q����.΃�C��c;��FHR���ߟP���6���*ڏ�
���¥��3}]F���4z$'+�������u�᪯N�$�����a��1w���`	��3�Vjh}���y��H�y���I���ۧ|��&����#yJ�z_�TGc�3�Z�����z�܆~����)�!iD�(���M<+A��R�!�.X��0	�s��;Fbհ����e��a�D�r)�\��ʦ��>�>��2��A����1`n�|�\jtj�o�b�2�9�o@�_��o��s:��@.�S�����rB��8����J3��@y(s��3�=�Emפ�O9�P7ވ���X3�Ei�:��*�.�`�-55�F�z֩V�?ͬJ��y���s�v&����9HGNv�����o�ؽ�\m=�]I�-� ^�BD�FØ�@Oq
d��͆���-E2H�,s�Q�L��jv�������˚���j_�Wꕋ(s�A��lۥIG�.рz&ֽ�2�ֈ%�ޥC��,ٝ2�+K�e
���A��7�.�IS1 B�����h��|@}=�z�Ӆ-��V�~��DvIX�wf�UG�KgL6��BLL���L�� ��d�dd�&`2����	hj!�A&����x��#@J��No#O䢤�w�$󭲃�{sY>w�"�Zs���ї�.�[U)V��V�'�T{	��۠�6�|g�!���>�_��ۛ�?�
��<������ۛ��+{�ƀw��꫊ x� ���yj��ې5)7�7Pݸ}���~��g{bW@Vp�D? �f���`f����q߿4a
����_��n֙�@��P��@B�����K�!����K���ʪ��y�Ą�4���=)r��@�s�o��j�3��B(o"v'f��M����0���\��p� ";�;��M��s�T ׿�@���T�?�&z�I.��<�Ǻ[��ɻ}^��SǤN�E����Z�S�>�D
���H�6U��E4�k��,����˺��v�q�o�u(<��Ƌ���v�4����s�_�[�P*�3�,i�]P&x0�wh�鴺Ǐ;�X*���0�_l���҂��Wl�,Z�)������B�ۘ�l�x�� �6:s��£$�W+��B0��V�_`u�*Rf*K���r�S���M�˦� ��۰�B� �����t�@�'����	#TZ�<�e��|~��GK���ě�Qr7��n��6�u�/U_��>����Px��[�_�^,�(B��6*(l�bE�}}�ʹ�u���lH��i���)���D�>;t���L3�lH1����cu�pA;�\Y�H�XfE>Ĭ������'׬�+�y�9u�h9K�Ts@�]�-�h=_e�$S���s$$���O���e�#�����_���1N�ua��.�'݇|����N�qƫ��x;͛U4�7���58@$ɳ�f��^v�����Ɏ�7R�kv{	FT�y�}-qPG����q����X��]�I:������0$��]��,z�l^1� �_�a��(�7����Q�ә�E�7�;�/^�,�ڢ0k�9&���K��	]$�)P��vgju;l�N#�-Կ��W��A���������<ܴGж���M��O��������QR��\@XLu�
r0z���lʴUu�ʿOa����	�'��F��;�gt*���7�
�!+R�+"�H�z��QE�� �d'2,�yX����B!�S`Ee�:����V� �oku1��[b���LP�����Rf���˘���I<�N���*�g��c�F?��a�����C(J��ߦ���Ӻ���^��\&��ar�\#�A�6����(���Q��|7�Y���T]Ua�䅻�7|�?��E�q�#2J��&�bRE�Z�r�MO	%_��½�k�\�肾H����	���ya3��m�9�����~ۓ��,_���D�nSP�ɤ3 �@�1_h#S&v{E�i�;��<&���үV���lC���M:3Y�i:Nc:�<�{f7��+[��&+6�kDE�VQČ�8v�V��&G�l���5K�g�˶t�ҷ��N!��"C�)����I�[}���2�s�7X�F��<kM���gK.���}V�����`(MyCn�g��K�x�D��^ � ��Cd��v��ǳ�4C�Iy��`��������i0zJ%���?l��"]1�2��{8�ē\;����3��O��kd��9�����|ǐZ����-܈�R�꼯?:��}R����sF������0�f��3,��o����	�F���s��c�P>�ī�x�3ͪ�@����נ�w$մ|ME���o�׃�,,�T������g�O*Y�0�RQ\}���mJ��Jۊ�#�1��7o*a� �H�?x�c��~���֒MAP����C��$��8�+.VlNܤ95��bb�0_<2�E�D^r�H
�v�N���%uK���Wz���
C~�-�_y�.V�oܣ�#�,���{����S�N=}�f�H4D]L;KL:^��Z��+��E����F�&���/xM m��i{��kM�1��Gf��h��r50I��F�c�(�+�����o��^
K�ob �-���g+��+:�6uF�Y�x|_,L�n���N�}�+����ҕl��o9Fr�\]�s&�ՙ����ݷF�[�"��5�m�V��U����(�)��V&�>f:�aO�Uʼ�7�ƕJ*��TW���]�wQ����3E�&ϙ,Xe�ꧩ�S��KP3����f�t/T�(���`+Y�`VO�
l����'���wC(u�tߙ��w�ɆWA9�W�p����"���_�]�ψ K��X��0@X��K��T�E6s�]�o�кεZ���p����"Z���*BDHE\CU��vi���P:l��54�A�Du�Y�e�a���O�="t�.��}�����:s8ؒ��ʷ@��~�e޲L,x���n�7}��2e���+Tw47��H�L�}���������w~��Fã��IT�g�)�%���"|X_�E˹�o�k�b%�:q@�~&X-���b� ���@�J�u��$k���*h`���1�%L��:rB5X0^ި!v���9y�^4g._���� ;����W��^������s��- U�	��r'^c9���
O5�s���:� 0��V�Z+�6N_��E[�]�xRţFPo���so��s$�x�N��1��������g�'�M:bм�:�����|��$�?�h,���]Xp�<h��J�z�"1��Uy�[����]vr�ϱ$j1X�S*VIX�d�<�bu�2=;ͳ6]���>�HW�P6�Z����b�;6�Yy��I���IJ���%�D���ߪ�'���XF]��y�e���ޅ�v>��Nx��4�J%��CZ�֚ߙ�0L�2i����aїV����N�̕{0`Ӻx����j�캁!�
��h|�r����-���dP(���9�L��M2��b�R�;k#ծ��A�z�U�z����dk�e/)w;N��o%��2���\���陴T��E��(�,8�w�9q�ʽ7��i�m&�~2~���P��t	A�F�b�2��y�a�dU@5�Q�S��q2�4�$N��E��3�(�J�g��\9]7�ILH#��;S�D�M��AE���T �6�*Q�
�i�ڕA��I�eT	Ժ��JR��*Ң!y[�����I�5�M#*��@����f�5�.�b�����w���J�;ś�z?4�p�2 ���)�1`(3%��땗'��b��j�%�B?WT{
N�hV1�*y�L.dZg���GED���3�ڶ1��%�v��	U�F�z�~���&jI�+����<"܆��ѿ��3�wA�%���֣�W)ă���ĉf��.��-A�GZl��'[C�Ix�y'̉KѴ�{6�5��'|pNMͳa`N, Tf�pY(9���@�zF���K�/�<�nbw�ez�ث�2��y/f����C���M&��{�R���<>˲l��,Y< ���δ�2iR�t��sxJ[$x���=�;�?�[�J0�~d����se�3�N��j�g�R�f�Q�̓`�N��?ӵ8��d.�PG�uC�!d]���LS#���D%C�ղ��Ι��ի�O��?dc@������N��{��s�2�hZZY	�g���v����Vu�i٪�A��n�^��xE3}�����}�����!3��T�YS�/&�Y3�J5�c�Cx��������(%�9��5j���?}R�zPB� ���B���:{�#��tvp����!5��B��aC�MA/��A[�/ep>Z�]~g���K?��;.��p�(���7LW������#�^��q�=u���S��	�Bd���/M���Z^���ӡ���yS�������W�m�Srk9扨���MO���N�5�N*<��yj�AB�z����kX����:�vj���}�>��B	����6g �DZy�x	�����%���莍��oa�Q�SL�䫫5��(]����X5:ʲ=M��V��4�BH�`/yHʌ`��PE�>EJƴ2��/�^x�o�!��C�?G�yU"o��(p�1�㳚�K1/�B�aZ��29^���V�vB@�ÒFu�?,� �[�;s"����|u ��`�tk�ʑ��XlxVHYEB    fa00    1d20��4�'S�h�e���_}g��:�2��}r�m��(���,q���=W�]�����;��ϱ��Yh�u[�Ap��XrC8�^��E_��/=u%�cT�~G�ʿW�gA\����Ib{��n��3σ8�>�������<��7���ē����R*�4��j�͐ =���V_Ag���/�
���C3���(��K���q������v��4؆L$���Ë���{KHH���+�^��	�����6��A�8�J);�V"+�^�JFK𴹉�Vq�q��0aӏ��kh�|Y��W/C�@B�}�OIz��'���?oP�7�A�H����c���V�	�Ɂ˃9�]�S�=3���,`�vo�����}P(i=[泴��.K^��f'������ݼKu�S�j�QV��IM�k8\�R��]��ODy8n۶��M[�L��A��R
�,�9A�Щ�����u�LX���a��Zr_ŷ3z�`�چSHB8a՜�jε��LU�/�oC�o'��RY[Y����n��%	9�V4�o����~6���A�^�&G����0�C��lø�F���5J��B ����^X��U�ۡ�����<��q<<�_ED�w�����n�]DF�A���on�f�捥hh����T��/vzSID��N3y��̯��a��U��_�{^���V%K���3]���'�ܡ[q��&�.��3��:�Ga����ݷXbn:�.��?]�����Iyn��L�����e`�w�u;�ԟ��~M��>N�Z̍�Vyq.K����?�5��v٨�>%+V��T��%}N!��Ѵ�ki]V����N԰��Zc����Y�%�"��dvW�Y�N�	j�Ǣ�� 4.�\ّ)�A�z?I�Yi�`�&�Pc�Hy�_쵎�O��\ƞ2@}vЖ7��FO��)a���0i�3����iw�w>3'[	�hJwmM\�؛���R0�/���i�y��/��Uxߙ�����};7�<h�l�]sD�W:��4�[�0������u����}�8�� x��nQ���Q�ܯy�����Ʌ5?cr�����9�:�kY� Zf���Ƕ��]����B�>?���qV�W�-a����׃�7��[��K�o"��/6zb��X���J
s�z�+�S�������na$��;�(A�H\�
:Z��T�gC ��X��7ǿ���3 �c�qq�Ӓ��.k!)�ța�v�f0Ga���a��1v�е��΀U������/��Ԣ�r_I[��T���6G��G�֤?�*@�v7��p"?})�C��\f+*v����`x����+��y#�&Їl.׏�����1�TK��i���ɻ�k"�Q���	႒+9�8��X���$�Ш�:��K�[Vc���W��[�\��+�R'R�I�e�(���uǖ���=�pb��w@ǽw>��&t��ժ�q0��-��t�2W�B [��j���QM	��d�i�F&�R�	����l�}�j�����ct�v} |,+?h#�c^P:�ڶ;!=P��	�\[�x����7?ę�/#s��"G��\�`#��f��g�Z�~��h[Ϛ$ �e�j��L�ɧ�ġ3���+���mӃ"���Ž�>s,����K��
Bn�� ��ה}��?��nynKeʁ��>ɿ���i�����a:�
�U�E,��TBF@�(s��W��M�x�#�".�|͘Kʱ��py"�wX^��Q�v?Z%����g��5X֑YNn>R���j)X�>���o �����Vh�Df$1U3RI����dg�=�Y����Ԗ��1�,YŶ9<�NB�y�3�����:���m�^-J��R3P�p��[%$��׈�<ǹ�k׏��ʣ��e�_�NoƤ�t�`���_�J�˛�i�#��	e�n��ў��0����M6��#E!$��2*�+7��@�OZ�i�� ���L�3�'Qt�D�_�����\����@�����ֻ�	=�����3x��S��f�+�B�;� ��d��*
��S//��+c<ҋՅ�D�f���p�@��(J(����BǼ�R�v��]K�Rz���B9��7��#,g��T���RL�>�ez[�䧱�z|�G��s�����$R�ҥ?�j�y��-M$�Jr�lEl�X���%�!0�K%f�7aV��yސq�c'���+�YW��5�J�JQ�^�2����J#c�K���T�:�6p냄Kqv6��G��O �Z%7�L�i�]�W2t#���H�l}���:������9���-�G��3����S�2�>N�Hg}�S�E2���R/�Vn}byK~��T��r@��.&�|�|紷~6%��es���d�2�Y�Oƻ���Zy����(,�?u}�bW ;ӻ��8�²eD�!�=d̺<]���֠��7��+ ���Ҁ8߱�1��`ģ�X���F��Ut�6?�Uʞkc�RĜT�.:��������-*b�8s��ԑcF�_XgKn�
�����o���_s` �C�_�T�1��	s)��4���Qpe	/�����6AN]�B���+�T���d�%�ׇ7Z<Q"�(3��F%~PVvq���MZ6(�N�u�<�M��0��:z�1��2�؆�}5ۆ��B��dlr�����݅p!���'��<�5c
��+b�roJ�U�MB�Jf�І���JH�Jf���<4���^����x���Ʃ<��Xl-�)ɲ<��384mW����٭��GzM (���7���e3���OX�?}_�At�a����Dg��Pb�t����킄8\_v����F�`9��
�~}�� b�2(�956z:}eK��"� ��oB�B���<�x�N�lj �"�^j� ��i8�뵘�]��4���*����(�۵�?�+��h(��u�X���1\JE�=���*;Sl��E�s\��O @�Rҟhj_`U/���֒�y�!�� �d1�Y���~��U��G:�dͿ�Ѝf3-��k*�1��dXU������+W�3�,�G�c��]C�JBZM��E�2�(�1��Я�1��佮�߃�h���q���W�B�0�b*?+����/Y#:K4�J�l�S�ق6f�����n�a6�;i�������
��WzR�t"嶡6��]0�>#�֔(ai��g���{�9��d�ӣ��4$H��&�w�����>N���C<v���9O��U�0ƵJe%І�X�e;���"	���G�v@���I�^g���r��DvY�l*��b.�&���Kn��;q��������ߑh�<�81��I-9L>���,&Qa�:Oi��C ޕ�$Y�Aq���GN����q,�U4A_��ibP��P�@���YR���5K^����@d������z�/s|�7)k��,�Go�����d�w�Lg䊈+\���_8���3�#��d(�	�n��E(�ޥ,�?����9`�Z�W<��%M�!O��8�<B]��N� �l:ݙ�7�N�=��g��vΟ�*�RA�ڍ��<�/�.��I
F��D�ő�Ɔi�Q@@����0�DӅ_S��z�e,�)E��K����KU����ޗ*htI�y%���V���Is�D̵5(�b��en'�(�r��62��wR��Q	¹����3����>�}�e;��(�7_��o9��H����~������P��z�2Ѡ��T�F�zO���OoO���t�9*�f6d�"�a�n;�X&�B �xd	 ͘9�1۩$ݲ��P՟9/�5��w;�o˗Ӆ�$��YX \5r�+ꔗ-�9 r�>�'����;T:��c7�#�w�X�9�/,߲Ut&�87����;��s�0A`$0a�[ӹ�q۟UW��l�A��bZ��{�S
�G��b4ܴ;�,χ7"�ԣ�sHTN"�����ӮV��!����m	aưѬ�4p�I�$m�Ω~�v�e���{k��R��� �ܧ�>���E��L��g�0���.(u��;�É.������`�]�+I$@�C%�Uj�o��D��5���#~�i��/�l���f��<.$zO򄂹4��XK|o!P��Vk%T�K�����Aѡ{���<ʍ�c�~��P��14��߲>`��EQ�-2�)����6�{������Z���F��B/�RA�s �6��}�L��%l��w�pZ�B�Sעo��tc+%[̗`u�Y�t�U$�d_�j�4|��#T�·a颸�r-�ͭ�zv�O�40����r��-�p�H9���!�'.�fD�c�i�3����~��p��]:#[��?>��k��~����8[F6)e�����Z|���M�(��K���7H
��>�ާ�:�9ȳ����.;�"�8d�n��:��6Iհ|��A��6~'�,f d�(%&��NDх�!�Y{ ��&x��_X�w2;�ć�����c|�jk��N��R�W�y�ΣG�rgd����Y��Ru�<#6��n���d5�D���}�to|tw��	dK����
�f��c��r���P�������(U�႗��/I�L�
����
��'��2��<�s(
u�����T�qab�^y���y"~H�Q��k	T�~L��Dt�+x���K�wz�4KT��Ў��Z�\�[m�.Ԯa�)CU1n@����'�ȭ���42�>�:l�O��Tl;�}�'m�ƴ��@B�8��4�}A'���C;:�L��hO�E*_,Yg����m�jAV~�v}Mj�<j"�f?�z�:h�Lᢸ#w_;�Y�E<��Y}�S���P�)�����D�������CLꁕZ��9�}�	����7
8WJ)�xئ+Clisk�V�b�-��?����,>�H\�
`�K�����[�)B`ﾐzJ%+�n���t��ț
��qy-\q��R��*�ˊ[���ɡf J`��AC 䜆��g���(>06؅��S���Њi�-��p�\�g�쳎DA�՛I��� ��U�+��H��*�C��-e���J���1g����Q����o��kjCܭ,��0|�+b��&v�&(q�t���� �����:5TK��͡�פ��T;f�XI���Փ{�<wN��F�Y���[p(g�O�-��:�����<=����p�3��Xʼ�c[��Ae�&X{��^��z�!M��e�P��qw�A���~��s=1/`��4+d �(H�)���@)'h�@
��|�zn���*9К�Ď�e������9Ӈ�� �:��t��$:$�;&��� ����p��!װh}B��jT[q��B��x	qp�Z*�3��`{�ӏ�t0bY����7$g�a�� Ai J˽b�[�a���hmS�a'��ˠt�i�bW�|'�[�<q���Y���7r��ȟ���"�f�H K<���}/��*�v�j��΃ߊ���$qc��䚡½�d�v=��z����9����M̦�t�_Ho:{)u��E�Ǔ��'�V��f����8+���Z�㰨����n�n�3moKۇv*_�,�	="1
�b7F�R��^6��B�d�ٛ�bO
|��_1��a7u�qs�֠�j�3�]5�
�? ��߄h�$C���9qI���!@�
O��c���F�I+!hLd��H)�������-ɬ�)�H\{
���[Q#1��;���-c̅P��YͰy��a�VC�/��_��|�S-v��c�]����l��d��"�al�#,�:=O��t�w�l"�*���W��]�M4��iﱿcYO�ɀ�u	B��?O�O��	�}����V�|�o��W{I��#RkIekj!Qp������@¼�=�t�}���7�Ǖ��ۘ�7a������r��ms�k����g�e��<��6�MY؋FÇ!~���i�O�oC�o?���5���<}^������ʌ����6�����4�^t�qlQ#���S,�B]�V�j�;� 	m��Ϻ>�؝#F�Q6Z�L��r^5��Ѥ� 5��`�t�-@��q��]|�PP���>�l��
�db/N$W�#�S#6��o�pl$�?j�����Z=�W��"���W���pR��wC&�*�d5P{?T4��62IL8�bVa�cy�A��e� ��8#�A9�:��5���<"\�	�s�^5����kC��S������d��y�a#(ԉAV�RW�ё����m���	}��_�@���[���� �5(�T&���	�hJ���mi���b/�A�?�����LAY����fӫ��T$�KY65��0am��� �u�D��Ґ-N���+����*g*Wg�E�Ǿ={���7���`��k�R ��45=��X���N���.oS�yƉ� ����i�H�<��ȴOX�ݿ��"� ۧ��q�d�|���dh�_�����1�����!
��A7�NʸBX*ʥ���Җ�g��FW�������q�z�Z������#^!�f"Ja�z`	۬b���xT���ccUF:�bW��'�J�o2�rzW�ԅ�V� 9Q�o����,w�:�v��!<YUX���!�I;挜��ڮy�B�f2���ȖDd��ʳ:z7vD�n�g�D��;o8wn��T�X��H��k�.�(�����}~ݭ0S���|b�s�e��z4�&�b�U$�?���
���ۯ��g���Nm��j��i���Kȶ8(�"UN��j������������k�'o�vR��S����a��lV14a�,I��,�$��(ǰS |�>�	攃]PP�3�^�^�	�H~�';�-Yw�p|e�*���%A�ȕTkU�3%f�q��T�cx�ha�@�6���K�ʧ�?��u�q��k
"/���AIi��!�ŕ;b~s) B�
"<���s�G��ki�gM*
�0B?X������q�E��b��J
f�U`��{�zc��W[h��9\a����(-��m�e��-����{�'x� ������.oB9[�i���gl�a��Ѹ(�a����0D��Q�dI<����%{���QQԙ���2��CI���D����Ũ*V��v�k���HE�`�d�zhpW���0��[���&z�Bܕ��-(+`ҷ6�7e�g��Ȩ��L=��D�,�u�A�d����?	}ؖ��;ۀ�>�*�݃���©�2���ā���~��5^�ץ۵Hõ�Z���v�j�/Q�H�dN���'��e��QԿb�0E���a�;���Lǌ�u'l,wMHS�e�l���i@�i���q��SO��ϠWy��oM�XlxVHYEB    fa00    1dd0
��o-eu
���i��ٺ]b u=ٶ�\쵖���B otu�
��( ��z9_��;�J,M�6zWu���"AB5Է{�	!b�c+��~��-���wx*��D.?s�!ײ�Vw�P�Px"ĜKY���u���iD�(@��?d��������OL����Ayl^�j{jL�8Wkzܸ�F�s��/����&/!/ɱ+g��.W@��cw��۝������VUM����e��cޯ���������������Ś!��MנaHf5���'�_�JwU�͖��;9M��j.��^W�9|f����>���b�C͆����InͺG^��|w��F�¤"E/�w0�:�B�Q��uTW���ODeV�8�86���Ho�E٪/�Q	���c�-l
�bE[nW_8�h�L��CR�#��D)�׺T[��:��2 �P���Н�Z�G�(?>m�����L�r�F�}�M�&��+wRn�7�?��.�{X�W�1�Ր�B�aV�\�SCd���u�����=U�ѹk�2��|-�0Fi�MT���`R<�ʘ1]�R�бҒ`�._�yMw02�t�m�t�C���7ct
�k��Q�!��C'��P�b�d�����@�;�\&�O烋d�J�^3.0
�j��kQO����J��.�`�ϼ��%�e�f��K�)&i�z|3W���� ���c�Z�d�7��Cc�c�R��#��9�p4��c�v#䅴��q�q��9p�6�ꍵIYW˩���Ke8/ͪu?��3ZaA��Sd����w��u�Q@�f9H�k~<��g�B;��	�\
\��;缠|�u$:���^굋���m�qM����c���!(k�)%�N�[3!�y-̆��}˔n����gE��b����h��pو�hg	_�AD�[�.4~������նk�����A�P�l\�6���ү��".�Ĩ�h�%+��L\9^��Ӆ�Ƃ}�hkg9'ŝ��uo���m��ڣe��Ci�q�cϏZ�h9R�e��o'�.U�'��NQ$�E<?�C^��M#���A~�@<)�y|^=�1�oT>��
�2a�����]�-{1{?יUi��!��_7F\�:��X�- {l�4M�M����l�����iD0���zA�z�y9�q!��Ytwz��[<�Sd0皚���C�њ�2�z�p[�B�߲�R[��[��LQ���O�?t�M]��:����&xF|7pO)}����޴�4�߅�ucl�-W�G&3RΝRKI�R��.�Cb
2È�����C�^���"����N��r?l��	@����p��T��}������<�Q��,
F�|�c1��0�
Nđ�����>��,�#%~��/QD8}xM^X6���oq ���M6?4�5x�"��
y��M�Z��,�7i�f'���J�P^QT;F���B�-���#7a����,}���O��!��O1��9���c"
�Ҽ��֒W
�M�?�� ݟ�s�畹��@��j��(��E����2��p,�����,9��V��
�A�X߬\H��T5�L����7�j>�A3X�b����k(�|�
rn_�����H��Ns�?���0;R�����Oħ��T���>���~N��5�[���p�����S�)�\�[���ql���6�E^k � �A�#+�Z�`�8Z�5Qd�׻x*�Ϟ��	�aO�o�K�A���8��N;����Y��G����L̏����"﾿��$�:f�x���������G(�|ڋ���CO�{h�OE�"J�â�}�2M�� '6��R��NL�3Ӷ5�Ҹ�W�h���k��=ʰ�'k��_��I�7�k[T���@�Z�8��W���)��7z3�W0��:�QJ���zE�:=�Ti_�55��v�Gr���Ôvl�y8!�M�W��|�� ��ր�&#�1�D�2�����g�*�����+w�ֺ��P�^��樟~Gަ��(�CǼ}=
h|�t*í��ӡ'*�.��m@��2?�y˼nIAt�[+I������8�KW�_�J?���o�.�����s��S��E�W.� ?�ut����B�������ٷ�*��]`����56�UU�ѡE�_�����u ���.{�A���,dGx��'�^-/Y$����sz��9����!�����M�N��K���}��)�]��j��t4�枆C�
wB����;�7�Z�x\�ϑm}�0n�Y�Vehg;��(�hOglG6�&�g(.�.Ȳ�9�
S����]y���5�K(4!�}���{�$G���i���ٕ-l������X"tI�i��K�_�{�����5q ����!�*���ߢ�U��S�(t��r� ��p#�i���`6�d�E��%\4	�dX¿k�����xm���9�/n�e�T��D{,�^��,���8
5�h��lJ
?pDݐid����UZ�Ӷ�츀��#�N+o�k��+�_-�9��U6��P��YXy���T�TXPsg�P�	9�ЅTح�N��qN$3%�!�6�

�򐾷
Ѩ���\�������������*��'7SDuZ�5�z�E�bE�n-�m^ǎbݹ�uX	�"ԍ�T��������4�����N�\\�x���:�q�s�!C)!<��=ڼ����Dh�+^�p�	��Ʀ=�uuc�ţ_�Jrѿ��\휝)��CV,�����]X�ٽ�(Y"2\���C(��<��`��>��;���yY��!=&0w."W���
�=������?�}Ƈ��*OШ)7!Ē��/�S��H-��q-�j4fH�j�ǰ�!����eˆ`3��`�� �ň#��ܲ�f���f������y{�Ӧj�bJێ~
`O�-���YE��߹�����W�9�i��u�~�* ��ʏ��錽�e���c	s���☎|ΔX[W%��Ӧ�������٦�����=8v���J���A�<a\�̸ZT#�v�r0�f��L�J��h�s4d�J����(��� UD����2��ZP�ȏ
2��!�*Vf���5`:��h�еr�d�q�k�Q�rG|���-�؏46�Xמ�u�������F|n���Y���� �⚬�%�$PvU����ߜ��ӫ��e�*a��x�@&�PR�sokf�k_�)�;C�F&�4�t�C��	鄉�n�r��c4���q���܈(�����l]����w�Z���؈SȽHm�.rP]�� =�yu�NQ1�|�cK�4;���l}m7�?��a�;l(�9�Z�+�/%���+����O���r������NZ
�7���[�`�ݞ�`��s��;}$M8��p=�L�
!w9X�+]���3&��GNd��mi��j�"+Y��]��Ja�=��6k �����W���<+δ"������!��P��z����2�����h}�D���q�S��V�����\�#	g�C�=�8�Q��T_�G���6#���1��Wn���?#� �A��uZž���l|.�6�X?8`}��ظe:�Y��w�N_���Ҙt �!x}-�w��J�TW�v��_�:�<!~#��F;�,n����6�1=qh{ч�;�*Ga�oGMy�@,`�>��ٻr��z-Kd��z�'�7N�2�D2����:!��P�wlV���a�����/]=Y�v55�nwNt˙)|�c?_f�PR�8��@J���?��0��8rq��0�P��^�H�ɧ�Ki�Q���;c̙O��ˆE.��}����k���Â�l���Jvu�e��2*���j|S��2u��\�!�-����� d�|H�~�P�J:&a���Ng��X��rEt˜F���MnC��3_b�4I��.d�1�'�P0���)@N�����}��q�PfC�x�f�������M&&�a懈;d��#:���:)H5j�
ɜ0mu��q�z�E��ڎ��Ԣ8���<�<V��?m�ߜ���K}���3.*+X��!��WoÓ�h�_������У#+ѓ't���P�Μ<�H�QՏD���][\>!W_YU�/s����sfԊ��w�{Wݦ�>d��c�i�:�ѱh7mz���l#|�m'`L�!׉b����g�͔4�\?�B�����º�
��c��(f��,d�~�=���A����Xk���5-^��B���d1��y˖�����	�0b�`a�&f�2?9Z��a�LG��v[~�;x�7ûx��K����k���Ua4��=��)a~�֤�$�Q\�e�A��_����=}@9�G���^}+O��TQg2����Wb`*�:��_��-���E"�Sٸ����q�2�\lҚ�8R�+�8f|�CQ��w�Uq�-������m��l�
�l�TG���mU�W��z�9j���\�F�jg �2V�7��4��L���D8 	Zye{��a��1����ǫJ�y��X�M��ć|�����S�$����'6�O�3�iZ+M`c�}WVu�?Ҷ�uɚI»K���?�>��^BoJF��1q�z���)1i,  `)f�O&������	�2�9�_.X#�>��)g�z��v��9*"2����oB2Yy44�?y.bd�,���'B�����oc��Պ|6T���ПZ�3�dh�\.��G�M+��u��\%%@X�ޠ���g��hb<P�Z%&=�n]�B��w.t�k����c�s�<Y���Ɂ#*��v�i{	'�E��_�Q���{b���5��/lY�.���Ǵ��T�Ao}m6BO�fz&|F7|���6�[�R%B�ŝ��?g���Ey�.���-�pH[���1i�߬/#�C0���G�Pl:^���{��|�W���\�:P%
���7W1��>*Uֆ g�
N�B;�&��
���7S��9gCA(�a��'���T��[M.�`=M��Ź/սϲIRPIDD!�r4w���-��
�O ��J��8����5�R.Arb����v(8p�h/C�Ge$�#��6�NUH<�-�8W�o�x��3�k���frG�K�H�P	�ߠە�����$������]i�J�f���v�E�?�Ǉ����`� ,G����J�sZC
tX>�2���M �M���Ѵ�L-?���z��C�djh��F�N�sw��`�ũ�	!ɚ@��	l�؅
>wY�����f��j~d�[��K�3��@z�&��"�\43p��!nv\�k��|)
'��E�<���¦<�N�)V@Q��|��F;�W�ࣂS�p��m=mҁ��Ô�L�w�N�y��EsSF�w�iS��9Gr�8��ٱ~H��* ����<\c<M�X�,�������=h��#��	�8\��ʴ$����h�� ����Z�����ˁ��V���>6�(���X�%���ڵ?�Q+=���e*��p��p>�4��{�E�=T&b��}��~.�ͤ((m�{���ci��ǅ��H����͕=f�(�t<�����I�T���m"�L`[F��hkre�*]��'����5����O7[tCl��0\0�/�̺����s��QO�#���bĎB�S�� ]
C�Z��%YH[X��RW�v�y��9�s2P�|���/��lу��Q��zL|��߮A�u#�Tm8�~*��aaJ�������yGK�A4����!�v��h�C�Ѿ�vri��B�w�UsР=p=v.g;��\`�>p����jX]c�!M��WV�b�'U�Q��+�#������d�0Y�մ���+T	�L˵Bz���L�E@m�		��.jV�W�W������8;G�ޯsA6���������~B_�9x�4���z����f:�c��rHD4���(h�x��G �|���p�jx,_�ɯ�-�=�O���>[󌭍_��RP����G�%�<2X�Je�2���7q�Q\焬�oO>��o�F�lvbfO��V���WS�����M	�9�S���W�	H�G[`r?��k��S:�/!��Tb���@����/�/ l�j4���Fz~���^����=�����/���!41��?��C[0�w�����7�<�>J�\��b�>��h26U��*�.����e�l��\�nwqE��� 5>�CC+l��`�nC�=ϻ�5���tVb�i���'6/_m�{����bƽ9��U���`𗿯��9�W�!�J�-~ƠW4�9�C���]����o�>����ժd�^d��Nh����y���6J�]�]t��6�N0��Fw���!1%s����]	-����ʐ~$���)AфNᷬ
i#WRH++ZN�54ɪ|#����#@��(���P���(c%��*��}?1�t\͏{S4��'�L���剆օ�����A'�gY<d*���^���u����U{����]��m�u������$��T���5�s�@��)�q���o�V lҡ�I8;�ӓ��d�bQj�tͼ��y��Bi��>��}i��r��\��	z	ˢ�޿�z�V �+Jĝ�f��1�x7��>�#��Ȭ���L�|��<L�!�y��l��=�%θ[1���R.q��I�j���tο.���TS��I��l�*U�8[^��:k
y�R�0��B�.ƺ��{��6K�Q�	E��0����4�_i~�+��+87�����(�����,��qp�[ы�2�ʊC�W7�Z�8�\�É0ص���K`8�nᶹ��@���d/����~;�
�Z:�
n�nN�ZIa�Ke��^�}�tz3�p`���;W���-R�����<���}�č�#�8]�s�bk�y%9m�r�O쵱i�R���U��p�Z�h�sf��(z;�G5���BScgs~U5DܮvSN
8�|*����|�^(���_Bj0����uqQa�c+��5H�}��]B/Qp*�$�fPE���僸�a���8�����7�ke3^���`����D��=Q.{�������8UY�;NS�����K��������x%22T�����7;����[��1xGmD�q��K)$��E�daTV�9��]^]�oj-��B���r0��Y���
�/�5�G| ��]폩�y���k�d��e����~���o��?����խ��Ģ&7UL�j©O�^�V;�� }�jł����P�HsO��S��v_�z��I{�̕�k4H!W�;�X��h#�*�-Vo���_�P��L�����"����4q-ֻ�՘hG�U����G����m�q�l�c�|�s8��G+�S��{�5����(#E��U�o-s@���`	�azL��� ��莙]�%�[y{r�pb*`��<ڸWQ�Gbά�ꐆ�=�b��UJ�ڒ�_f1=&:��%6���"�A�]�㒩�TU���E�9��Ql���RQ��Zpj��w�҇�8b @���ʏ0J�`�XlxVHYEB    cc25    17c0 �J(����<Ӫ�a����>��S|��w�P����6'��tg�q��6\b�r�T�%�F��Qa������١��=	Mfh���1;�-�k���\����p�S���>P�� .h�t��{jv�Mzib������K�sl"
�+u�y��+�r�[F�'ˎx�|�%X�>�Q�#��[gvX�Oʬ�?�J�栀�w#Ĵq�k�H+��{3���U�Cs)�/�����ήKy�	�o6LM�����vv��8j�$WMr�L�@���Tr]lS�	;Q	K}?ذ�K �G^Tڅ@��[�#��(M��ʣ�i��h�(f�E �>�N�m&^��b��{J4�x��[�c?󒤶6,q*��d���JU��������0�����Ş5�ԣs�=�YX�r�λ24(Y�BZQ)�نS������+�[�l}���W����N�����u�0��h�7]@�%�L_^fH�	�EKˈDX�#P�IoE�e���&X���
i�ȤŠ�+��Z�_4ݸl7	R#�8瓡�*8YL���r��Ց73��,h��e�s��|�-�~�봁�G����b�ի�|R�a;�ZJ��$HU�ꩾt*��ZF@b& W�����P��G�@<;ͬv
#�5�v :z�� 0�	P^J�S�����$�N��b��[�q��KV#�Q ���X�Ǌ`�,�P��K��ǡ�道(���v,�b4k��I��пϢW �Λ*�}�/;������L�*M.�K� Ƥ�n9u�^��x�*���SDg��H��T]��7v�h�q��D@YPk�?LۼK�a=�󼚋��_T2BD?A$m��ӳ�SP�s��G��ߊ��	��	B�}]eM�2p0-�Bȋ,��p������A������s��x;�YX:�R=y�n���Ѷ}�>�,�c<��M��������1r/M�a $݂��wȖ��"�"��?��͐���w��:���)_��C��<���,���
.kdnS� uR�/��Xb���!���.q���cȽB�s00��kkc[�UP�����WХ�et���e�]��aͮ�[�b#N�y6~�)�D��:>��
�O��������}��6���5H�P�j�� d� ��k��ۼוE��Z'�v�[��X�F`6]�Jga�jU1�&Q������'�|1�$�J�6 7���hKJ�R��\؁xoֺ�-$#�5��y�`����݉��K����_"�tM%�w�Ŧ7{wm%_-�d��¯C�b��y�Hק�f�0����l2����|%�Y#�KZ���q�nt
�󢅜Y�R����h,��@ӣ�����ۗ�T���TʶR�>�B�1�˨� ��8����'�X�c�M�= 	�BK���PxZ ߈KQٱYVKg�T}ף%�)�{�y���?L�����U`�(�l?֚�ɭx�3��Q�Qd��i:
��%�1,:��aX �ɷ�A~Ȏސ��;�6~���|�᳔�L�/�WF��9�ҴHi��^�hWrn��{��GO�^ Q�`^<�v��KCá�g�.o1|���=(6�����M��(Ϡ�,�>�]*���
�
���.�����tv���M�f
%�^f��Ͽc��Ά-?�*�~E���=R�΃1�A���6`�g�
�8R�_��8'�]�����t��"�d���h�e�d$�0��H�b�]�ig^�����V�N-Lt�rߞյ���Υ'&ԏU-}a�䅗~���.k��B�P��&Uu{�x%/��l��8	���1��x�hu%�ḳ|iR�l��˖�7"]Sm:}�@���1��*�B%�_VC��>uk�L�+ܮ�g���]W�����f&ޒi�&Q��3g<�T���*���"2���k#��u	j�g-�q�A��ijD��tjA���+�d3�Tp/�7��3��0xh�j�k(��d��3m��9���:���F�g����wjeū�5,�\xRĕ�P����y��|%�{*��C*׋���<3I0���ȶ�JԆ(�j��􁭞{�]�=����"���L=�(�m��2[��+e�w�}I�o��㘄���"w&�_��(P�@{8�2r<����^d[�Jv��`<�G<��%�$^�-�}�o�cV�֢�S�0&}3��Ȇ7�B�s��C��4V�T|2t��٘w���O5,L���p��ѵ؊0�ּ��T��Y	��f�W� ��=��(^5� .��!�Ut#������Cu��@�xØ���@�C�k'�û��kj��lD�r|�$��V����N�4�85���\ ,u��h*M0u����f�vW+Q�9-��Tn*'�a�q�o&(�>�����x���HS;v{!܆�%>�!��ȸ����^�4\���(p�S4���S�	 �W����L�1�Z$Uj'��{޳E�'C)i�l���Sx��dʤ�-��;��x��S����<������V�N$��~һ��>���[��ɼ�{��#��p�� ĂK�������`eqw�T �l�A�{��U��w�S�E
�����w<�f���d�(�M�
P����v�uq-�����=�fH.H��c��d���}��c%#��py����"F���^�݌�>o�E+�������Y��
耤�e�2@Ȗ/p�h�ۂֆ\ϧ��J>�y�+sI���X@��o��+b]k'+8���y�<��A�o&�f�D��5?��C_4u䠦_)=�@��L�И<(�����#��ZxE?I~7��;ѓ�	���J��䷭u����篗a��u�}���%�#��Pk��E� e�2@Θ$�~�R���q[��1�>�6u��j%]N �BܭF�[=TM�!sV�!�R-�uv:����������g�և0�\|gny&�����q��:a��֨g����1<_ywRt9C�ؤ����-��!_W#�=�7��c����<WS]"<���L�3�*��7��IX���;b��b���IK�$���?���R�.õ�5��D���iu��I���~��h��$�!��:(S�㡛�� A�&|�Y��]3��\�73� ��:k�-��*Щ�<&�_C"fK���O�깊*$M�n8'-HZ!�R#s�pV��=���M�<Ŏ��6C$k@Z�����X� {ݵmB�����ԼV�^�v��x�?_�A�	�_��l��yM��[��1٢1�F�R�3�ҏ&�U+zF��� �;ɀB�$�[�F��Yp��ԥ/��X�2�\v��6��|�|@S�!�&�E���WR.L�8%fgn�4W��߲�<�C�1E�*�������8� � L�1�R���r�%��i��EtF��c��f�#�����S[�4���ǥjCXv9.���l�B�l�oc�mǠ���"ew�b��%I6��[��Bzv����0��r^�6�/�wЈN4T�$��l�����.-r��`��W�X�����U希P��*��`���)�%��o��������[#� �qE�H�Ư�ЉQqТH����h>[�PANeGv&��e�Y	|����,�h�V�`��o��*��l;/���@礠����9~�޴k���Ve��2��̣�Xƣn^�8rǮs���J��~'�����<�'i���sd�]O����g��� `j�#�CYOgݻ=ˉ� ��0��$A�u��?���3o��3z��M�Ӏ
>������<��N�L����~�=�u?�<�^O��?�u�d�������+"F�jF��Fg��2}D� �@�A �O�Oҏ1c��R�}P��N�/�>���Ӌ�2K��V[a�@�4}��»v����]���RS��Z�'�2����7=�F�+���U�d��/í��=�pK$���x�\���4� ���%K>IZ�w���C�L�U^�ܺ/Z�ͺ�� {@�ޅ�<k�m��D���P���SJ�Ѱ��s�g�5l���k�`5�,}ϰ�|p�rEvĽ�fR�uG�"
(;�|��3gސ�v��&F�f�.��У$��*���L�;��,?�����(x�(�[9ў`�Ϣ0���ڸ!�}+ ���o(O��diM}��K���Q\vt�n��o��AЃ$����'��K�Ul�o�菣�<���-��MǍe�ue��W���J�����B�ee��]���oFq��1 �(+3��y0g	R��ZM'�g���.�� 7�����`H��L���U�s�Ь�wz*V�1�ƽ�s��ͷ�q]��в	'p�}��=�i��o�-=�;��J�S�A���1U�h��OK{���d!Ue�H����7`C�J	`щ�qgߣ:�E)�i@N��E0��n���"���5���>�$l
������uh����n$�?,��_�z�M�j5o�]�+C��b���d)+�r��1�~�����k��z���WE�"ӻ�h�³k�:|�?Üu����~�����T/��d�t!wN�r�>��+����X�E���Y�A=��zVp�i�����s�s)��(9��&l��(������9*�s7��tp^�~�Ѵq�[������d߈'�"}	��=FN��&k�3�����mlEn��-�g\m ���U[�P%q	���`3��)1r��;Z��,ݩ�%����A��I,�� �������Zu�33���^�H�t��^qc`{`/VabU���놮=ΰ�Tw��ΰ��T,b�&����**����.�<0��[�����P�u�;���yھz.���?�D�l���,�*�ր��3���O}��mW=���2&��(�
ܥ�r���`��$%�l���H:�J�-5ҘFHO���a�NgO M���t�wi�iX���>��x�m����h�Rf�+-�����ٜ���X�j�=��$F��1�.fه9'ų]R�.���F���;Ƙ���W3`m�w�l?����ߗ5,��^Ԭ��>�;@;>W,�A�̆���a���՘N�Β���'�',ʾH<owH��y${�����)|��N���S:�g�f`ڑ�t��
��0�C�m5~g%Dk�����\xw��
��Kwӷ����f�?[_	�� Ո2C`�D�?�;Sul1��&r�ܖyL���Z����;�t{���@5�	`Rڡ�����9Ѿ*<�/�y��h}U��c�ԍ�_��)�	�v[�>�� q8(4��$���~��ڴ��X˴M�6�2���5+�WxSS�E��q6��=#��H�Q:=��}R�o�'
�h�̬���"��}�2�f&*�I\�`ShQ�����=&�V���v���Au싐��Ojb1.Y�����E�<�/�����A��:�D�A'����:w�	M3��i�%�8
����࿲1��u���a��1��6Wq%�dU%e]3�m�V�B5���8>|qr�PV��H�u_���yr)��q^6,d�����Q��-�5�p���K���euO�U~8!��x0Ѷ�2#��� BG��h���k�)ʔg���֎���?.T�ƻ�F�x��	�l�o�s3z�H ~"����1 �-��n��v<i���*K#�V��4$��s[��~���`��>@�,r|"]�*
ֿ��[�5P���U>~fI�g,	�I>���k����Y�����6��J?!\�!���:�br��j����^���p>c��$�\�@oR�����!Q�w��˗�|�z�hg��n�0�|5Oa������
�݂Rt�y=t�7��ЙiVOi����[�̀�Y���P�my*)����)	�ga��&����g|�zQ۷�����9ZgD]Q�1��lk/k?>���1C�
B�}�<�!�@�,/w�����7����T �.��6�;�!�@�ߝ*