XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����$�]�}�Ix�%ә��nI�Rcf>q!gn�Z����|T�J����N[��%I�2+f��/���*|��s�h�V�$�j;;�k���
jM_�(����{`F��8�<h��Qz�ۼz�y
�gl�qNVz�ϥ/m�vQ;���K�M�^�949,���j���'��
I�\#���Q?R���̌Q�n�?�n�pN��@T:�	�l�5�,[&>O^0���=h�D�Dr���l��{~J!�>'�����l-�Bڙ��/����ɏ	�bOK0���8}�M6�a�~]y�m���G��K$�:?FX�W�ֲ�"A�F�)���g�+�(8엉:�4�ؕ���.��=�c��>w�d��� OU����c�|��%���C[�a|�l�[㇜t�ߋU�&�O�M^��~�.{�����y;l�G !ҽ[��4��\�
��i����֎���"P�a�T�x� wޛq��e�7z��(s��A������l}	$���{D��{	#7��}Uy��S%_)OE�����6f�Q�sԋwc����~f�w'R؟E����(:�&o���g�7*�P����Eȶ�R9>��r�+� ��<Fë�c�I�wY�R/�!o���hH5F=�o^��Z����K���ǎ��i>�O��5Q�@xN�Q|jFF����9�fj6~e
�o���;��;p�&���YN�	��v�$g��n�vp�!�g��㈐�t:���5��F�Ȯ�8y!� ���v��.�tXlxVHYEB    1a5b     890XA&�5l�͒��V&�Ƅ����)��sTֲ�T���ħ@��f%������R�V����%x���X���2�2[U���V���P5
�g��,��|,:p��j����o�̄�M&�����k��oe�Zp�,���*,NW��{�Y�X�w`^W�&I�I+`���r��~|���,�Bxgϝ�J�/���R�+�n(��w���`�On���ػ�]F�g����'��)�)��������D�[ਡn��2���c�s�`����XB�/�57��oMG]����/>4Ŕi����u�Գl�+��L�E�7�7C����L�e
���ջ>���E@�v]H��;,rd�z�qچ*��Y���V'ߨ���Hڗe�ۧ��&�="����\��\��p�|8���ۡ�@��O��MR�<�1*��9jv���J��R?o�������%�b%שw��-C���`�5хjDd���q�� ��l+ĸ�H�(c��W��n<>���R��7o(͑�&�V<�JD�þYs�K<?�Πt./ϓd���x�I=�,w*��.��2G��vMh�@+��¶!>dW"1�;�K��R�,�$�Ǡ-�y0�����ⵖ���K��CGB����0��l.�b�wo��%��i��Ep��R�	R���z"}��i���s�aw��D�r5!�H��.�,�!9���T�mԛ{������0Y��m�7pQ�v��O)c^�����2;*�V8���2	E�r�oI�vX�"W���$q$���m��#~��7��
�l�a��^߶P�'7�(i�%'��W7�Ѕ����)З�=j�?�{�忠�h�����UT�ԩ��w+�^1=��h&a�I��R�M`|���	�a�駖�}G܂�4&�4\ތJM��A�_����M�T�yF͓*�iI�D�M��\��@��ԝ�Үz�qBM�q������ZI!�ٌ�h�E����z�p
8&q�M�-����S�I�*q�MM̈́/���/���+��.�P'3y���0�fZA+K0=�d��PS�x�	z��i�|��oVj-+�ǀ����!h��+}�^����VY$�B1�츊����>���_X֩rBͫL&Ĉ4��/������C=��#F�����48�å�f�Lǂ�#���ך)u��� Hbw�e�i���9��6K�\�#�b�i�'I1�f�'	��W���IC���؎	��-��깴r��VdFƲ�ǭ�A�Z���Ý�8��u����q���6V��H�\a���%�`�
+�TC�&m@�Mc#[{����O�C�M~1���s�P�~���W=�7�� �1MS�N��P�F�)B�O�Б�`�x;Eb!�]���K݋��qZ����i���I`�%��Vc&�����99a��Y�q�+`��LT'ݶd�_Y���2m�SE�ћ	2Z)08]޾�f�j��Fa��N>o�8sܫ��2���iV��)����_
�砼�1OȽ�|�N�cK�ػI��D������mO
�̼��w6�K)�3���j����a�=�<�k�o��ѣj�>Ye�I=cGz��y���ηw�$�*S�����5-eTfIW�nĚ#U/,q��h��of�
�1�Q��zI���NM���_�q�;�<��I���L=�/�<1������H>"�F����B��o|ath�d��������IM^��Cz��g�G@��3�S.�>��׃}'|&�u�D*�����L����0/;�,O�?Q&���;���&4-�e�}Ȕ�b)�4�!�e�tb�f"jr���PB%�d�BN@��
 �/��D>T��+=~#�a��T�I��K�p�F��
'�	|as���sA�7ZWw�i�f�ē����!�({��*�����G���t*���3M�;��)�[J|��E��\F2�	�0��x4v�9Q����o-L2�x�z��α�v��w��kc�*j��iA( �.6Y�oسG ��5gB�yl�$4$���.���&E��x�HR( N	)�V���i�7�{���lx�h�Ga��$��E�b���>���1B��&f�|��C|���{��p�̃�ͼV�W8�5,Mk1�x��A��}2G�MK���	�9��|h�{����@�g/�: