XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����"��7�h跛��y�l��AI����!ތ��ȳ��K�	Z�c�nR-�`���K�Ͻ��t���0�yP�ư|���tυ ij��XT����;��x��z��f�og��Qn�:q#��O�������Am^�IY�^�A+����Zv��#�~��j�eI-}�A,=��k�>��b�k�����E�%\O�Z�	Ĕ�Sm�%(����&��68e&X�G����ij:E�9"$;�)�m��������O���`5.����\%�:R�Iݳ&��ap�GqP2r�D��7� ׾�P�r�k�?����9�z�]W��	��p��0��am�W`�*�B��S��]��^�r�Uk�4%k�g��6�D��&B�⸟&�Z�(tj�l�,�I�{�gu\��a막�My�J���W=H���'���(�_�`�E����g�W�����}�3"�����f�7-��:\K���cA�2͢�Qwv�����w)�G�.�'�&�i���_�i�G�tF��>9v\Ud�b���i�:9�|�A�3z�j���9����MT�6��_4D��>īlo�8���ŠLl�6�㬻�.�� �&3��U�����_M�X����I��tFV����Rh?���,ȸF��ZG`�����H���MC��dE�yR���.�1L���f�Y��'��xp"��Zo,��6�jR��G���\i?�EX�h���R-X�IL"���@�c�@Δ@�L�KՒ���x�K{��XlxVHYEB    2cfc     c80j�=YX��z��Ťه1���3�/���EK���(��^Ӥ�䗔��=1�ېvkV��pVA�$gn��OGY�Uچ��SA���ھ^U�b;���n�^�2L��hh!j�(Ҋ��F�V_)���wj�5�7��f��]:\`'� �`�ds��A4�5�K�(���{L#gl��>6gl�����:���Sf;\��N�ՠ[D�rn��Z�A�z%��pj���8Ժ�EU�H5�E�T܆Y��$���"<�A�~�����Y��Y�Y�ٻ�0�(T�NX���n�{'6�f��g3�̉��+F��Po,m�"��9���e)�kX�T����N�Xa�
FZH��qу��p6f��������g��t�V��i4����O�'�J�e�)�^)w0�܀N?�|"JU㲣^{p�^{>��mL��}hQ��ך��hv�~gQ��M ������ndw��n��m�@Dw�!$�����5 ;�ђ�2�n)9�ZMS��#f�n+�@��`����@O�{�x���86�?�U!�����g�@���E�q����k���)93��H��z�����k&�}!WÒr ]
�L�I��ոU��l�?-ƍ�3!+�г���йf����X�G��'.�0x]�&����&�@�ܕf}~ED>���WgN[�Y6��v� �-����C��hB�!�q���?�p_��OB-�0��u˒�TuDyfs�/���������I�d�_/$�S�m]ڴ�B7AV�Mͯ('	v�J]��[��#�����Rǟ�Z#��&�	z�-���8��_�d޿�{��l𠈥_)PՖ�]-h�g�˯��������J
j�[E��[v����X��6����,<�i�&_�i�y���)��"�=����$}�����f�?�C�R�0���S�s~�M�BW��g9}�b��O,��Z�[E�x���J�/B�����D�%=Fj6�Ϲ�8��v����=h���3�unu����q\=M�8����ד��-�f[(�0�_r
��$Ʒ�fI���M�9�-�h�����2����ڟ�A,V�T��0|�x��}�1z�H|c�f��B�v�����>7��v��D-��t�w���*�?�bOj��k�y��ϯ��0cc^��n����iCK��>��l!��8Yr�����O@��F��Y�z]hWG4L��9�Hd�=�X�M���e���%^^�×m��J �w� ������Icv�Y�i]X��I	���u��[u��ۋL�j�g���g4j��Q���rا!���`{(h3�,�y{����1�,I'ήw)M�5j� ��8l��R��tU��������)��Xx�-��������v�]y�����,N!~D��S�=%+���^��aE�o�9J����K.*���-��Z�~�O&E��޵��X�O�I���1�{	�S3 7S����*�)�wk�W�(S
���\�v˲��O5��Яȷ�UUܰ���?��v��u�p�V�g�Z��I�� ��lj79Q��2W�`��B��'���%Z�g�c�xԟ<v(�iȡǙ��δ0�&��l�O<A"fN���{�?�v�j�ȗ����#z�&$_��;Ap�
���M3 �5�f��iGA�x�#	�%��v�h�m�؟� \ �K�(]G4V[ ���гF�e"%bW���.��u	O�̿�ֻ��*��<i�c�b�	T��ץ�_�y�c.I��r-vǹ]H�w	�Bw�Fe/�r���g�P2md���h�
X���X0W<�(bJ;��Oh:��\O*D[AD�I�vaY����MNm�&A\�<�������D�����.�1A��blʥ<VSJ��E�'�g�;/�pOlj��lM����,���ݶ��k���W�f+�_(0�w�4���'v���iGk���e������Suz[�s9V�F�b����R�|>�\�c�*/@h�5u�n���YӞ�l\|c�
�M��Jj!(_�p���ܘ>�
��n+��y��O[��ۄ�>�8�}1f���8*�0 �l,A;�m�V��̵f�vX����,��&K��I�-?{�!������eLdzt���I�������=��H���'G "�#�*����"�\ �o��˦�]ݫ�C.�(*�y_ZePM�d/���+~�3��
������@Ѳ/ey)�%��ޤ�i�]��}_�D�o�1AH�Ɩ�û�WcV.T97HT6�"�Gk����d"~�W�[-@���R�[���/��Ko��i}	2 	��,U�'p��99��e&����6~f�W!�g��}�9�9�KT̡Z���m/��Z��Y']Ks��*�(�F�qD�=i8��t�X��xE����?�s�[�׿�I���E�-���ҕգ��.�>����c%��ٯ�D����zȐ����bp��O��[tzl�.IY��,�����=��ݖ3�ڴ�uG43��j�V�^�#S�D�Y���g�}t��^��A�s�r$CH���;�_�P;(J��h��j]�l��ja�C#�s�P������Ƽ�y
Cvva1c2=W���vT�&@��H4	?}据��Ln)�ܝb���Aj�QZ@/8G�#?,��pRb�����:
�j.SG��Q����{.c�<gF���j����"GG'�A�m��I5�̖H��G��K�"����o�p���Rw�0��&]Y��:��?	�6�b�t���x�����T��|��i�������v�m�4A��m&�l�7�a����D��ƌJ@l2��q�;菻87D�U3��!`
�dh8U~�ig�H�f�����9?i��-����*�<�;'���#����&��)�D =���4?BP���l�X.��vꜘ�0S�E��������S��y:j�+���A��j?�N����&aZ��=�!���-Yz`6ή�gm# �)���_���3�5q/�]��4�ޖ��.��"^g�	-��!��=n�l�!,>��Z0�H�x_Xt�kw�#��k=[����Qٲa�Ն8��������:P�~�~&o��1���6S��+Z!g���y�}r����d�s�-��E��S�4�'��#m���Q	P#�	�~5�L�i��DԪ����