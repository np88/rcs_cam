XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��r��2�z���L�,%�?]r��m/g/�xV�u���cL� ^�V����'���`��;d|��pr^d�l,�/?��y��E�%�~��݌��U
	i�Qc�#� 8=}I��
s�u��WjN�߿L�E�,�l�?�Rr��J�-��D@V��	���|�0�k���]�Y�☦F��J�K�N8�^o�(���(kż�ԑ�:�3�@��B4����ǰP�'kt{b���E���Zf;;���FSmzvѸeEi���nF���x�M
rZ9�ãBP�|�-�`8�1�B�1��Dn_Uг����)�N~��b�঺T Wǯ�M�f����u=:4�xF��JcfmYF[!μ~�mL>�s�Fp������WԹ����D�����~�>�I�,ąI�q*׎)F���Y*/��� _ƙP6����:~J���&�����]�+=}^o�&�Y���}#:y8ذ�4a��}7�9lYTЗn(~'x�t(I yb��6S�hN�^jAH;��lA���:�V�n�PG�.GhJ�w��̹�P�+A�� �v�2�Ge���U8��֌���3O��'���$�qG���Iu�)�D� pWpP�\���j�V��"��)��T<J{HdzϿlIZ0l����d����B��B����WѢf��U�i)����Sp��?k�+���їT O(�F$X½f#��&����
E�J���$�_*]�-s�	�.����Mr���䊒4��!�e��Ӵ!��$`�XlxVHYEB    29da     af0���@*��ow-�\�0����ɳ��[�chuQ���7:�-qw�6H�8 ����s	׫H�4#���{r��q���ɱ؄ ��R�DP��[�ݰ:�ґ���Wck>�qJi�������E"D?_�[�G-����̈VTG��CbѤ3����y� ��)hG��fp#
�h�-����qu~�W��~����;L�����IBp�~���Ml�+)�����ۢ�Z�ܿx�*��� �n��Х�&,)�W'SWy�|�Q޵�)
��1w
���	GP�J��ߪ �O�����6�SP��]���tX]ݖO��A  W�`� ��@���i��8��KUHM6%���)��% �^0�x�����j�'B��5�g>S(�xP�JWKQ_V����S �B��sOmU��j<��;81�35��	M����Y�f&f�Aҟ���Pw] �02���\�� �%�s�p��,�Yn2H��]r{��/?c[�qV�ifF�5]] ���j~v��|	zq��l�-���5:t��/�;m�Z�T-+���j�@�J�H{�ʹ��/�y�i!�=�.C3mV��֕�t�Z����������ߣ�Y�Ð�L|��p�����*�e�ˤ����,@o%�Vl�ܕk�īW-�d��r��B�`
���JD<��v5��?c��~ 7���� ��yJOj�П`�@�{��|�+�z��lqQOJ�D����z��GPȫ�_9髰��'�t�f�O�s������ }X>\O������k�9`1 Z�+ �S�u�[l��qeR�۾�Z��y�ܣ=#�j��@���R��=��%�ɢgme��2�X-kZ5�w���]���ͥ�Uԟ�p�nqZ��)�C�Z�#�%��
!dG�b)"�7��b��c��g��QR϶�W����4�	�P��·�������9�%�<�
�O����*� ��T�?Q��\V�]~���ZV0>��g��A݈�#C~��x8N��Kl|�|�:�ABf�	�u��倮�gTݽ��k�)�~�|4S��}- ��
�$&�Y���#�x8Ű���
�GQ��3kuF������C�-Jv��͌OVi�#��L�(z uk�!2�uZFxKY�/���������J����ǧnM��,�vk�>�����U���}��D;���c7�_n�L�k�#d�FN�*��(,憸3 r�Oy�m5�)I�l��o�ԓ���š�	
�7�-y���.(�_*Bf|C��(=����b���`�#i�ŋG9�m5bbC3�4��)7�*�E�~.A���b@�(	�~[����́)X]>���/�.�q�I�+�L�N�)�W�څ�h]9��4Ƥ�����[T�]�~�ۦ�����w7ܝA���[�8U��Д�,g�W�P]gO �C1b�y9���Bt N'�V�F��PK�R�6թrbBf�\q2�tp۔��M�H�w\�O|���(��S��G�u�[����{��rb�c-���	!+�^
��`�Gg.ѹ��4� lk0���b�g��s�4
��"W�����'���!$	��x6/ٻ��V��&,��y���_�Ag/��qF�QM?-�Hǎޕ4Fҝ��G�
]%r$��1�HP����"���>G��1�IaQ����kq��cU\J���8Y��[D�t7+�>����8��%38���TKB��H4UV�O9r���Eݦ�"!�C�po���n"�(e���bH�:���&�Z����~D]@��J��2,��d�m}�����)���%�(�+e]�LY�ڽ�f;���V<y���q�,��7$�ՠ� R,6}��v���Q�y������F���ɱT�+RK��� �@fr�C ��tvl���_��P%�ѸR���!�$��(�|=����68ɭN�;o(�'�>���[[�
�a�}�u< �m�TeXG�8���˹�U�f�ۉU�sa�v�Ko9]�9���o���o& ̣d薉�I�Ӻ��;�!ģ%w�o��P%>�L�;�l�v�}:֪��gJZ}:�}�!�2�I�JGA%IdA�w�Z�'�#���XtJ��R �"I4Ug�ke`Lc�m�vi+/!��z�H�|���:~C�u`�=�?K�4	(Y�(�8�VSx��4��cܷU�������O�/XA	��[�%H�Rh���<.�׼`9c\T�T�oS��&��hj�1�AE9��|V��"*�����:���� �YQ��[��B�]U����������>uCN�dPH��q���=o�s3�//�?�o���и���"8~��w�\�3��W�;��Ӿt�w#�����N{��&$�6�|�K�n�������r,���ӄKV�T9���H��f.�GI�?����)f����G�x甹�'�A��$
��O�}"�)�eZI�f����U�pN�E]�sv���޻���Ue2����.~x��<Ou�&�����R3���13f��vБ�Ǵa�ʟ~���23PW�m�W��P���x��)�p�����W͎��t�쀶��8��� �j�s/t����Cwف8�rUq]�%s�o?'T9$Rħ�ༀ��|�d���J^�,laj�0�GkZ���k⼔���bD��
�rL����1��d�vm����N7����F�kv�i�~�4429R�H���b)�@��F�~������+�|����9����ʡth�X�0	ʔ�@%�v����3��e�3iH�]�b��#n�F�H���