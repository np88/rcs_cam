XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��b���ǫ�"�	pUg�=!�=4�9h�2'�8��f��[-�:u0�JO�[m��G��R�e-�˼"��]��R ���#�N4�4=���q+���d�մ�� ��<!w�ܺ��Q �X�LD���)�, �v��/���b��t[�%�m�y�v����`��j��"��6u;�#�S`	�(�3�O�~��ɩ,�̌����Pr�,�P$����V���e^3oj�ӣ������i�u֔iM,W�Q���2�?6�V�Ùk|�9�鼔8�		]J�E���O1��C���H\�w}.�Y
}X"����n��r��8�\�K.{�7z<#װD�?/�X��'!�����ei�w��vw��o�Y]F�V���l)�>����ڀ�C}e�e��g��1"��_v�.�����tI9�8d��s����1��,����,^g3���2jRZr�v}a���H�j	�$���C=�Om�f��ntf����0�BL庶����X�˪p����,3�
���7�5�[$�`Mi�|M.�|����4��t�`4�yzpq0�u����q�
ٵQ}\�L����S���z<�'��2��q-(N�5��jY�-�0i�������&�q��H(�>��Y/PJ�9ʉ����~�F�����<E�!�f2�&�x���N�Ep�w��_�T��36@5-��r;��\���@C�[���;��B�"���;�%�f�Cl�v�3ȋ�vk-�J2F�e�Bk(���F=��q�	�_¶'Q����}>7]Y-XlxVHYEB    125b     760��A^s�[ϲwG&����ܙ���62'�r��)����[w�h�M�b�s2AJ���xq���0:L�-*e"��tD��1�ף�W�ǲO�ыB��H���J�#'<�;��P���4	�g�3��	�֬����9��+Z0!f�vy�9q��b0��;٨����d����3��4��d?B�1�[���;d-�i�9r�g5�~ڜ:�����7|t�BI��+E�Du�7�n����"��oR��A�c���T�+�UQ��{��n�\^D�;N���WP�tC?5��ʣe n qB���mu4�HX�B�}AVغP�^�$Q�2�q�� +�8k9$ş٣*VJK/����[덿,W����I&�����+��}����(s��J��Skեܯ��7�leL��]w�i!���P&r�w�o�#Z��$ګW�	��-����]/���ɿ�Ny�]�zYu=��?��.�{+G�����x̙��1xDߌ,|�;n�MÙkP(9�l��V'�'��aʤ��c�0�G�l�h�����7p(G�^ ��V�=0z�Z���������r�[����z)}���+؝v"F��c�35k���?<�u ��� S��pka�N+6/�+<��Y!l5)	%uK�Wp_w@�5�m�'(
��l��� Է:���Ů3 �2ܞ<}fZT�K�.K�N�<wG�=�
S��D@J
���z2= �ٯ���%�?g�X�=3��{��(��0��d`<4�rG n��W�m�c�9��8nZs����QjG�gVs+�m���5�e�(�T�QBE�X��Ϛ�i��-�N�YV��F�}b��^� X�r��K�߉����R}�&w����ޠ���R�!$�s@=QS�w3a�v�
�� X��������>ꌾ!�.��32����jU�,鈵K�7��Cc`�r��H`%0gn�e+���0�^�+�����5�X�3��y����#H��3��/R\�2�.��"Ү&�,�u2¨s�|t���<`��,в���FEך&�o��>M�ğ~�D�q]�K-G#�B����V����}��A,S';܉�����N|�J�~���*�6K��E�Wɤ�Q��n�X���VT(?l+�{�5����+-��������q5�j�7�}���FhzlS��2I�����X��"�w(�x��7B�����e�7��ܲ�� b�m�߃�n>�R��
�[��{d
C�T�cD�ɗu(Pq�PڶQ/��vgހ�����=͟��B�
舘I�K5ušg�E\݉8K?�����_��C���..ڹ�C�I&�`��Vw�*�ԡ�-�k����Σa�W"7��d��5��{|���C�%lIEgBR'������<����p=0{�/f�@���?�K-��r{C��f�Q@�Ȓ��qm
����K+ʻ�cdm�@�\�d#�j�q�2p�����oD�֡PG�FsVG��Y,0Um<{�r��K���e'<�w�%���������� ��,�o&�W�h)���(���^ c�ؒڀ\�W���6��l@��� }��"/�q�9�D䦇D�F���{d�(�kI�ǜ+C�NTp�:���>��"�[�[.�Q��<�z�m��_�|h��m�<� �B>v�NV���'��U���h�Ts����pϊ7���ިTW��O�"��̓����^�c\�5Mg!b�ΐm*t����K�]b\��I�?76��=���[��G87�eQU8�h�2���}K�Ȣ(-=�}o���j^7��YJy�B0SK��6������抐7�{V7y�(�$����d��4Y�K�f�C���m���x�v2Qdu+ �[0�8���,%l�5