XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���>�!�>t6i��Z���C@��Ԡ}fk�!.�Iat~����Ӷ��t�%0�$�LK%����K��osז�gq�B��yQUİ�4 Q��[��N4���}��t���,ؿѝ���3�J2�]g$2mV���lH1��
0)#���$b~;�E=��؀�?)��q�����;8�}��b��SD�C$�N'�C3�%F,w	��$��i]ɾSk�2CǙn��W�_�/�9Z�7�?��a�C���k�<�"��&�_'m�����G���a���	�C��1%q�*,��SH #�R���p��\������(6��h-��!�#�g��l�0����!#/	a �U�3�m"Yb,�E�e�*�kR1��r���-�9��.��π��g�OG� �nn�������V��r�Brb�d}V�5�����F�������� ���n�+����̏�H�`W4Z�Mӻ^H�pb*����%��Z��	���մlȣ�8��¡�*5�=:���,������"#u|�K�ϰ>�um��t#[��1�ɵ,����f*]=iԉd���TZ���'cO������^p���v�&P�ŃpAT��b�?�vb^�m&wn��ۀM"+t*�����$qtq)qo*����^��7!
�P�b�s!��Y#������G���u#*�E�L}�KR�v��Q����a�6��h�j�:�~��1�s�F�2B8����?~7>�����镶��}�q��Z��YUu���9�ד	YSWXlxVHYEB    c6d9    25d0�e@S��4HB�^�K� ���ꁋrd�N���2�&���qV����v�ī�6��Dw�f�h���%��&� �
�Q�l�B�Za5�xG��ן���������K��������Xfnf�d���I��yԾX�_|~�6�|�Ӯ,�{R/O63�q��Sw�\�t���ۡ;Vf����"8�8G@�=����
ڸL�t5��$V1B�~���t��u@�{Ѐ5k໩+�S�I�R��7��5C��v�����|��s���D��!L�7,���l��8_@��1���JJ�m��߼�V&�),a�F�^<j/恳��͍=�Q���+f��������
��\q	e{�ٴYZ:�(fN���]���B��
�Z�t�)�N"����/O���f;��1��tX�-+��Cvs)�	�,�3� Pp�bKT�R�=Y����.!	K{y�Q5�#`|���C�oP��I���_��ƊJ��	+R���A�5��D�p#�B�#O�N3$j_�>Q1q*X��v�>�`j���h�+yDCr8��m��ܥ#M��V=�����P��]<��;�Nf��eE쯖�
X�����;�Û6�ս�a~�p�.�i����$O|n�؏�?��ȜI�~���o���NZ� �������`��� /=�B�#Hs�������0H�M��N�"z�{v�V Ǥ�K�i�W!��� ���转oFw�+�=J�\���u�7?��7Q�>�Yyq"9,,�	F�������_�������M�G�Ua�r�W��)�P{��z23�	��ѣZ����$G9�2��wXb6bd�ؓ4��n � d�U�;F��.a��H�X�y�D?[�;�N�1�(����5�"�%�t���0(�436hF �ܓ+ ?��s�#�<�j,�2L6��\%�=���	�W��[zH�قW�*�z���0�w�ȘT�n�L(��t�{e��f�4$��8uǚo�c,����Q�[
��+#�4��0(�M9��3�����I�M�Ȟ�X4���~��[�q8�:�iе���Lx3���CN��~ l@u�i7��+'�H���> �C�ND*�Ӿ��P��5��J��3+o3�o���O�
�&M'H)�m*�N�_,?N��<4ڸ39��'��GҏG�߁��^�/�pʜ�W&��`�c�{��7+�pv0�^��'ߑ�I������b$p���^.��A{��)���������[�mb�^�A`��N�ecaa�E.QqP0O�H`Mj��2�7Z��g��F֦/�t��*����#Uf�pߤ�������40��<a#�o,C~KӡfP�F/Wһ$���u��'Rx��ir��Ec�� 6'
��ÆG)�pi~dU���4F@s)4"H����.�ה��3�l,�X�Z�����X���M�e���c���C'����͎�a{Z{�ݣ��?�X�10u>�u�o��Z�� W�6�����l���_RH��R�5CӑjZ�>ԭ�`���n�1��"�*=[��C�?��m���5됲��c�]�Y�\���o%˔z�g���:Dx�=G����Us�*C����{����yw!��k������.�s��I�}�A�Ъ�O�V����
�[}Y!�sC)�$��>}Fyu�9�	O@�8N2:�ߪw�	�n���VĖ�x*�����&�u����e,J٢[a��*��y�( �R�^��ײw��Ϯ� �H��7��s[����#2���'�Z��ް�sF�����;�_�L�ou�U�4X�V��Ｍ�\K�D j���n��2�BN����Ά�j}�pF��Κ#3��b7R����OVmY�C,�`������l#2�p�
�"%`���2�}�½���`eS��Q�_�kU�h���|c��8)���^<Z{��z��E�������R�u�c՞c.�A�����D&���k���-nO�@dփ{r�{8�{~���21O���og�������c{��yt<P��f����IZ9<:���YH���͋�"J��ނ�=����1Q�S:!��z���WdG�O���*��y4�����=��;E�
O���4��1RF(�J��S�·�n��Lw�}��^{����=g��t�
�%A�h�戺�͛O�w�3���Dt�7�\A�:Jc\k5�w%�dU����x#���D���Oz�h*w���X�I&Ց��s�~(���MMs�[хٿ;:H��x��V����V��/��%�N�VSW���\���Ō����N3e!�j�	��B�O�z#'!ѰVX�t>״hA|�?��ӕ��T����� g�D���]iƭ��-�Iy~fL���}�ӝ�Ό��*����\%h�>�"�;d]Z8~�*o��,l���ω{_��_��lv�8^
�@����Ym�*�֣����V��Վ�<��R��о�i/��J�:~q��ybB�<��_D~��������{��=�
n]��scP	8<eE/ֽ��ݏ�� ��糽��\@�N�O�E��I�Y���t���6*�n�P;c5�X�5t,'+1t�J���B�ʔ�Cu�6g���CC�,[^΂!��T��r��w3ѹt�=�-��75� �k��n)�o�jw[ �u��[�<�WՑ���}�$���TJ��F��C�N�Tؐ��H+��Ｈ�r�A�Tl��ڨ��s�b������Z5�k���y{L}'��;^PD7/4X����C'�)`̝p���@�3FP�/>��|(��A�F�Џ�W�Sx�犘ݨ��`���G�mL?�۹;�^� F�@�E�z#���u����|#Y�y���?�9�Y����Iko��]p��w��W�N��.���s�*�2�v�B����$;ፙ�T��vAfH��yɣa�M�4������D��`|��c���uR(?@:��G��Nf�:���J ��v��9wy�_2r����}ѐ��EY,yOm���~�z/���fR���V�����[%�p��%�!�a.��tY�W�7���@�EMv��Q�Ӵ����1��װ�ȉ��4E#���v�d�@vFd$_@����mǗ�#�r�w��٨L�n�(n ���@'%��jO��{1�Ք�6�`���Ț_�q�{�.������_�Գލ][���1

�(D�2�dE�͝0��< �Gm^fo�=�����A�j���n�,Z+��hu5?��u��D@*��!ͻU7)5j�x�����c鍌쿴�m�͵��p�n�XM)h�`>χi;B��I�lʠ�t�х/]�X���C�V��6f�)¸A�4����m�,?�Q���x�� '�@������� 3Ս8F(Zb����tM�Ȭ���ͳ�;=<$�ӆ�(V�����:�n��ֶa���4�i�M}���|��C��)���b9c3��Cf�|��#�����.�G|�D�N��a�c/�65�=����������R��OV�bl�<hu��X�ZH�� �W_O�WZOy�ѹ�c�_>�_Q�2�-]����M;��!��,O�Î����J��}qD�
����h��15���y��T�v�c�Ͷ)�P�QU���L��$Zb��NH�v��ϑt����cC�ם8a���_����$�J�|�ado)���`�p�\|�����^��^�e��,y�i^�ip%<�OR5:,[���mNv�P5Z����equ�Z�y�Q�T'���Id,/q}$Q�����x'��^
�_��N����-�&�b��
�qwe>�ޤ�LK�[@�Aٚ^�K�!G���X��o�*[@)Q���^����<��jkPY(��X0@Z:��c�$�8W�W퐑��DVPW}�cx����֥����a;:���I�1��v��gO�)���.�d?�?�z(M5�i�)�ٴ����(\h��&����n�X��D1�����ˡ�7�K Hʧ[��͵��"s�6_\(�1�9�_�Gpؾ�7iQG�͓C�I��s�`����=;_�-L�mC	�DX�|��Z��j� ��"��4UgXu����	�"��Jk�µ� �Xo��[��ʷJ���p��� u'�.�2a��5н�(cY
��¹ɂ؅
QQ%q�i���DF����R����ܯ������\?c���S<�9�2w�+��1 ����)O�ǽ�8���׮�������L���J�(	|�}�xV���!}��Bh�T%�-��=?9.��]�(�	��5���_�Ə��@���Ϣ��Z�;�c��J:�k�����_�4������1��w��s����B�-Q������8t�Z���
ߎ6�R(c�J2�ex��DK�*l=����:�F]�S��*��/X"DjRmo��cp�(rC\�#66}��28A��u޴	K� !�u�bVY׏ny�>B��VC�A|�a�b�b ϲ3T�'J�?Og�!Hn����Os�� {c)�)��LT�Y)�$lH݀ܵ�y;��lVk�V�%F낒���p�B׌+�3{gܢ�N�������k�}w��6S~kxla��t#��P��a�`'�y�s��W�D������χ&��&߈R��煊�1H�4מ@�ėq���	~�c��f2N���?$Y�Χ]�,�p��e�� )�����bH^��X�Ӿ�BФy�!��i�e�C�b(�ĥ�^U|v�J��������{�Xw�8G��	��,�/��i�Y���r��-�8ᗶv��)uj��,�¨!�*ne������Ӧ���!�ל[�%N�|��\��YD����27�ƁJ\�ՉW�u�/��*umt�ڼj��2�9X��c8��#�s5ko>p�jip���I�;��㪻�hOP���ʉ����0�wd����ek-����FV���G��Qh������:��_Q�o`��^@"��d���r�6!o{A4@��G*Z�l�O��6i�^��n9�����L�x༽k�?���B<�2� �3��o	���a��S8ҋ��/-79<��Yo����=A�U�����E�0~V�s���n~.C��i��ֳZI�WƼ�����v�Bu�@�#n�Z�$��V�����2�4{<P��N�.ZT�y,��E�,��Q��v'm�e�噘R���Ոn0`�,�j���>H��<�
����v����Y�5и��_�ہ�dW��6w�l
0Ϸ�, �=����fT�����LdB��j���h):=�'՘¾@A�,G�rZ��A:�s�;�X9%ӱʜ-H�g^��|�绒�j��$��>�[(Ƭ�m�}���o�IAM59�x��kM%K��)�����D3�\�Pv@ܪ�CGQ��?�
+���.��Nv��}�[�+��5�ɉM׆!��폸���oP�(\�_1�G�R�� }=��@�Eq��`3�Z/]���}�R+d-fF�"�/�%�Kv~$d �#gK��U�1��=;hJ�AM��=�d�G��L�G%{��{j\"P?�)K��������ߙw\<ں����mj%�S�w�J�1t�m�Tp-k�t�)!ȳ�j +C�=4[��J*��-���5=�M�����(��x_�Ӆ;2��A���M��Jt������8>�ĉO�!T�Ӗ��J�;fEώ�D(;�4@�G��V	�܅���yX�"\�|�P^Gz�&5�9�V�B��K!�� �3Z���U�ֈ��uq�*����Q�S�f����&�QR��`yR�i��Eq�J����1˩��3�-�r��3I�P?�b>6u�5� �x&��BQ ��A�<�c%�#����<D���߰>g��P��Ā9}YVV#r�ID�-5X:���Ŷ�	�S��f�}���>���&C��X��@�x�	M2���dI��pp�l0�E
�1*�I'�E14vH�9X>�CdH��k�X0xt*2���k����E��4,���B]�Y��������ZԖ$�"0��8F0����IH	Ŕ�P�=~�禿g�KNjbL��ξ�HQK봗v�v��ʣ`�u�1M"0C!��Ƀ|�"6���B4U�}�$9�wCg��[�k�SiK��������q^�:�҅�Z��|fx��y�9���m�W�soW-������e�tP��K��GY���n�
2�����OL�;h��8�l4��`����lvX�f�@+�MCn�e&'�F9��l,�z��Z�,�(ޠ��ކ��o�C9W/H �.[�>Y��Qn�Y���P:�1$��c��8���+QЯ��b���Eװ&X���W�1�l�Mm�qA����}�!���7S>HC]f�������8����I���Ջ/��g7�xSV����n�1@��Ԉ�h�H���v>s�+��It�5t=�k��Ҟ�7q��������zO:�|��J%�ү����?��R^!�����Ԙ8���Ƃ1����E��mt�C=Y�m����V �
�
��w]5Pq�#R}���@_q��n�_����!�o��K�T�\��N��w�/��gH*S]�*]�[ژ�ד�>���S�ҧ���B�B0�
��@V�C3�I2bDn�Z;�T16h
U��w{f�pf�^�⫩��,d���I���<�d\�8H�#����We�e:����[zH6*p��-��]5�������Ż,T�V�Ig���N~��3x�K���$��p�->ޥ��zX��\&U_�d�!���vB%�fm䀲yut塍:��"�+m�i��I?���S���[�{�3���ȒF.<>d%��G`���>�xH�x�}���7�!�����ٴ��)7ݣ��d���P����D�)	����Z�*�3�I ,f^#̵�\]e8�kFZ-�&F�9�i�������EZ�k�^��'fF<��@v�Tg��p���ې�`� o4��?"-l��GH��K�lҳ~�"��E�D��ǜ�ܑ���F�{7��Ԣ�D7��of>�b7[�T*(s�.��%1�
�,X�<։�D~9Wn,!����M���Vr��CL��s4�J����C�h�|)�G?��0,r�)|�$�,Ae��8���X�J�T���s��N�F�e7N�����f3����ä@y����W[�ox��K2B�{e*d�_1z�V(��P�/�sP͏J��d.x�~������Dj,�\q�-��¹	�����2��G��_�k+>媸KQ����>�T/�w�%�:���P�����q�< �����6p�G��ذ$9�?��;7y!�E4�Y�ZQ���. �r4�J�
��;8�J=�>��H�`��e)�_��?yC���[�J�P�L3�5���N���!���}���;�n3gd�v�&�����vЀɴ#Ll�d��]��eL
�\�n�"i{��^b ��d�Xn�>>7��y��x~���q-E�~9Y�:)2<�ӡ�����,����:�+�2�[<n
�i������,�`G�i�W$��vx^�w���1�JP�XD�2�@{�����C. �nv�N\�TV���X�&Q�r���^��(>xRA��Nۨٗ=�fiJ9����AX�E�E�( ����O��"�,��6�lXX�N�G��IN?%��d�	�ȘM�Nu��Z�u
��M�R�D����GM�JS�y֪J��Ѷ�Љ�i�x��$���i�1��M�FGxg��)Q��$�9Z6{�=�~����0��o���M��8o�b�0�ҩ�k���e=U7�!�6�����)�n[�����h��H %/`�{���Dԫ��8��$�!��iHL ��1����rk��`�w��T�cJ���Q�y؄��Iz��N���U�c �Oܕ�z��)p�[>k<S�hzG-�q��=ݾ�����J�j�w�l��;�Q�v"�AVJ�KdE8)^�=i�raC��S��S�<�x;��v���i$�y1mR�<ku" ����F��ܶ�Z�~ ��9����=I\���">�N��SK�ti�략	�P*���R%�K{���5`<��
�"��+���k[�r Mک�(L��d(��!V�M��_��L���F�E답HQWW���󄳻<�c"��b�4c����K��$�ӵ��0�o]���sD�K�؍ga��q���M��	�I-�sQ�a��)�b��d�����0#�*w-�/('��F���wV�B�)dv�)�����q<����.��s$���l{�:�@��@��?L���Y/����;�J�M��[��p����W.��_��4�	�����=W�G`l�]TvR@��3:6�gmЕő�|�e�P���2����w{B�XG����V�;�䰭 +�j[+{H��n�lԡ����ZA��4 ��&�3ckaf�3��ra?pG@Gt��V��P�����a��#�|;m���8!i�1���x�H���E�Ih�(�jj�j�������������0%�7��o����bڲ��',��N��ՠu��E>��d|ngі�@���+�a��rA����W=����y��r���i�����i�� Q�(��Ŀ��Mr'GR��a�l;@i~wO�!���3
zͼ~ؗ*���C;X�J��'��������G)�P���e�~��ɷc���Q�imo��|���{���S�F�B�� ��ዴA4�`��m��j�`�1jܼ�>%�6����B��_ TG��_BxQ�lT&�
�[�k0��[�K�:5oݗ�r�S _K5m�5���a���.��x17{���՜�R�Y�~] Jm�j$%�^߅&�M��,��Sǅ�{lRg��O�ҹ�}]�Ӡ�� +޷��?-�P�����1�-�E�$N`��c(��%�kv>�� 0S��6[�,gA����b:�o�2{�G��Ku0 *��Z�N�,e8��3X��7޺�up��b�!���ܬE�<f�Ͼ��>z�^dV��%U=���.7���ds'A}x��r(e��nsݻ=�ǲ�f�c��;�(�=�9�3�G�%�셨б�u$.�͖��P1�?+-��ܪ�Z|���
�D�7���,0Hk*F
~p�;��gP��1�.
�P�^aj#Km)Z+�j�(He\�o�;��-L���5H�=9e�F�L��Wf07'S���bԶJ<vl�V�f�t��1&&����d�p��a��z�8ڂ`?݉�{��I���b�)Vzlch�`�p�#��-�s�z��Xn���T���K�]-�CK/B��͒;�g���.�z�d�ՉY3�8h�y#�;�eNŅ�D(��Q�Ӭ��+V`?����I�s�&�n��B����A�Eɒ�RJ�DX4o�������$k?�A��[���"�4]��	j����S�х3ǋPPM	��>H�=3�y��\0R������˓���({$)?jj:֮ �16s0Gf*��oc�B� -�\�j���F�������]W�r	�n��k$�>[�!5[v������S��