XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����hHƶ��~;�,�E�C���}���		��ܳ=��Ҷ�-��s�#->BA�^��mw��f9��v9��]�QE��9�Y[����ZR��TZ����}/ Jk)&�c��vs�����O�B����@�6�n�����;nI��~B����3,}J�ٯ+�8Y^^�TNmu�������yQ�P���Q�m	�}���C�F }L����6]Y��6*�p�B�b��'�W��QC����r,;���3��zӱ���_�=z��=�xm��/�sS�L"�N'���j��,a34h��0>�8Rԣ�Ih�p���*o��D!/�A�`�H�Dn��"i��5��8�+�l>Pi8萼���	�ڀ�*��B��c�D�6�u��ە�3&iߛ��P_-���?���9+��R�+�m�C����.��K���?�H�A��s�Wx�"o�l�����f���9��G�e����������e����ò�	�Y��U�.B{Q~(@S�V+���M{��d?��$�������� �V潻gJV�Q����zf`\n'
ª:	��s���&�,�d+� }�����K!s�ZF2Ar�s�R���������)º�!���i?mr� m-�562�֯4��Y�坹�o��U{��j#e�GJ��̊wOI���e��-q�ߵ�v-hP�1��
���焼�5{�����G�OJ�h�s"�p�	��;�K(ņ���X�Ô֮��m��^Jf��L��vH5XlxVHYEB    3b6c     e50'��5�5����!�w�����8�,[��g�>�J��p�r�5^{n/+d��=�*٤pr�%��:��3�[#�A�[��꨾�D� '�tL�i9N� �d�Cy�C�<�FY��uCQ ӊ�_�W�sh��8׭/I�h��'N��+̽yZ4�����f���:@F�h]i�]�T�G^P4����
��F�r_�'��
Mt�qw-to�h(�%0���g�P�ے��7�r�ۃ\캺��J!�@�~:p�@Q���2]�l�y�pjxۙ�%��F���Xl���V��@�)/�f5ٯ��rv�%�7�����a �B�z'.\^c�{ET����2*�B�'x,4�7n5�D��x�����[��L3���C��v�e��Vy8�;��J�zE��%�RN,��h6>�k�,%Zč^7��>*0�1�*�[6�D�q+"�Q˰[�9@��
���M�7���F��:]�)�K�!,l�|�	`�T=�߆N���ų��ȝ�Ét��Y�5�b��o�7$�/�~�rb^�U�;���}��	к��6li���y�m��394fP�GIE+?(K��CȂ�"q�>m&r䦥5�Y��0�fq�<��Ŏ%pv0�sfQ�����8K��z�&2ǀ�o��a���p��t&K��nz��fr9M��ة�<�{"p�o�*)��Uc[� �H�'�( ÷[��tb&d���\��Rخ��s��Y1.���M���~�f���Uq�I坤�z'���vg5� 6('�����f�F /f�%�ue5Z��$�WG,��n�����|��&�qs����u+m�fn�����IJ�ս	�p8R�q�f��L�VDT][�����]�g�DG�y�GRUeE,���Z�iλ���1��!X�O]�CЫس*eQ�������p/�KgFaG��X�w�B5�a1,$��$H� #��{V�V����WW�"��F�;��88$f/��d(罏�K�n��f��b��?S2H��s�tf�ϡՔ̀����,�ѝ��mڠ����.���YSU�^�J�[��@źm~2XӿR�|5����1�ٺ̧�Q,Ȭ�D�c�O��Wa�+��x0��R�㟝��lra;�=�	''�������M�+]zX�C��mZ���$�J�L�t�� ����@��+}�B;�cĪ��ީ�MtU��6������z�i�D�u�10�xi#�,/�?��I�*70y��N�a*q�o�C�
ȝ���y�9��n�%^�;��N?0��'o�~`5{&v�Ц�[w��v�}���Sق̰�ė�pId��yV�3X!{߉r��X��#�1���Ӽ�	��b�10��̇HA��"S?<��y����]�?,���흣�>��,볷Kr�RB�d��
���٣��E`.[��i��6g�H�\�l_��G=5�N����5hv����ؕ�����F*0bq��y^��N��=��L#U/,�H�#A
~�����b��M�R��\\�M�9���H�fe����OU���^��C+�.��E/���C9��X��CǴo�-��*�n����!�����2#o���:!cv�8}�|�?��U\A����� �˗��,G�{���>x�9�A�MU�W7��ƥ�%���U5C�1Kq��0����B/�����yܝ��&��U��"���%wli$>DW]����PCZ_�v�a`����0�J����bܭCV
������r)�3�Psfn!ׂ)�y}p3��M8�m
O�uk�3�#���0�$�"�wJ��Tbt�V��9Q_�ee���v���x��3��Sq&ͨL�qq��#�<O�y�K�WO�1��|����v��a���n�7c�`�b`�N�����-�(�`���FK�
���Bj	v����'(�Y��,��QC++��}
���f��T��QsK����W�����v-RS߮��k���{�z{�.�80�T3�If������G�;���D4�8t�@܃nF����j#�����+�Hz�x�K�L�^�n�qn3ZTnT�,��d0�}R<"�p�̌��ߪ2ļ:�C�4�8�N��;�m�4$(�[>�Je���Ws�{��ov$���O$T+����^��J�	#�R�b"E(����c����V�)�g��]�I�q=��K~+D	�#lwڭ*"%ҥ��9)>���rM�\�X���I��,B=�ה��U����cdo���
Y	��RVdL�y9-Y��8z��!?į�}����/֑�y�f��4�%�����K�g��8��9Τ-��ȹ�ӱ�h/�3�F��c��d:���"/ҝ�[��nE<�����N�7q��[��=�)�l]�z�����3��a}В�oS��N3�N�.�]����矁����?��`�5��:}����.wF�k���R�źv�KP��)������N��S;�A[i�9��*����
���P��:�Й�!�rJ�R�&�=�w�F/�s�Z��IU�� �Wl1���6��Oª|{�A��L�q��p}�U��M��G�g�J�o7�/;�pKP7�9{����!���5�hH2�.74�`\7�����V������Iݧ�"�v��Ha*? �����d���M���I�lc�j�Bi�r�D,�؉kf-�u[Ҝs*��Q藊�c!r�<��o2��ґO��lg��Y��.E����$�[��-Ԭ����c��&�ce�'���j��?��� 5xq���o����_�����D���3�ps���m���"�����I��O�l�z�<T���I��EW�<��2~��q]�Ed���7��r�*[������˃;�%Y�*����5�Iٞ���.��\����=?����Jν,�kk@Ok�9H|�FOp��u�Hl�����i]�Sf�V~��ϟ�E8�jx�u&9��:�&x��f�z��V��L{����7�H>0�����̍zs� ���83����9���������;ƓT4��ն���%�5S���NH�lvaЏ%܈�"���sH�jJ�t���;���Fi�t��-wUA~�$=�
rV�6r ǰF@b�XL�ε�d���xի�$ri�qc������&fp���!�|�Fګuq�����J�;�xo��Mǩ�ӏ��(����;���?�1u9�����'2�R޽���I`�[�0q��j�D�t�Q�8��j�#�9尡�l�K�ÀR�� n�^�=�������-��)_�MTjSI�+tu�q�D0���G�>����^I�:�<����t�ί�r�����!����w$�����]TW�� �M��q@� mNln�_��gc'��u[�Z�Gf�|�M��y髼�tcjx���� V�/��sK[��h[�?��P��S���?�
��i:p�����o�g}O�:|zڃ��7w�c���4�i?���^2��>H�G�6�x�|ll��P%�찌�b
<Q��׀�2��?C����� l�!鴮�P��[N�+��!G�mM�R�� g,��!�D}����и���sͶO�����4#���ׇ�v|l�ߊ�T�v��n,]|�"�Q���[7~��x�