XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����I��+lX���Ty�.��^v�}�s����7�IҘ�y�|eܾ�������?���9������y��!^UUZX�ͻc͟c-��^ZZC)Ir^7A��|�Px�3|b|ڸ/��J��
�Γ������	kq&	�N3���(/"B���-�+={�h�eg��|�v�Mw��!̈j���Vm��}�${%�,�PR�����5�W��i�J�P|��a�X����-W� �����c'
�I�@��Z�;��>����RA����#p�@�8���d�G���%QNɄ
,>%2P�iyx�q˅�(T@��a�N��Y��o�z�/&�Pg+ש���Q
� �Iִ�}5��-;���v%5�鿌4�N��6v��$3'�,�z�ϾC��txs�s�wr���N��d� ��NOMw�1�fZ�����njn��:-۞�p��b3�D�z��d:z^�>� W��;���7��/��:��G`Ϲ���V��� !��?�M�ke�̹��\����1D���H��R�,���k��HZ�h:1fj�'Ʈ�Y���jw)�xy����Q,�s��N}+�u��L�g�kaw�aj�c��J]n�m�=� ���,P�%D駓e���W�@�����l`����o����*fEH�b�yh��*6%?#I���G��&��Zh���۬1UN���
&��_���1'=�p<A�T�����~A`˛�AIJx�m�q���ُz���!��_�n�9XlxVHYEB    4cfe     dc0��"Lި����FJgv,zf5 M,n_��"wl�'�.:F�ޘ���d,��B*���?)����HY��Ѱ�7��S?�� �N����r@l���W��l���Q�#��b3�h^.+�s�y,I��4Ż.��]rk;urr��;��!���?�N����m�����K��I�X��"�[m�O*i˶�=����s�յaE� �p�+� �Ba�4�L{(����Zi�ޮ8�:��0Vm�H�&�������Pqصf�ql0� >3�aa�ң,�mH��"�;���V��=��v&��~��4���m?>&�䣟��凒����{�>n�*��Q�q%���ֶ�ٴ0���x����uN����x���a�(�c�x�?�����4V���F�Cj�K@�WM�*������ߟ�j���Y�%~WI~�%�י{m��o;Ad��5��)����Z#π�[�(݋m�	�[a^Hv�fe����W�ŵl�c�1�ٵ�˥����)b"���bO����ȁ[��S*"�u���ʪ�� _��ũ'�y��ބ?���:ێ�)�dq�l�V�27;�I�ɀb5����;�#|�.�fDA�0��rTW���C�J�t� DH�P�! �g9�+iJoK���|}�� F�waW��c�@�b��D��. zi枮��0~ў�PXz��*:¬��eY���y�H�ɰF\�$B�����4j�X�y�̐�8���Ϥ��s~i#��n��e`����8������0[�;��ŽAig�.�����A�ũ�����W�z�9*�����6~�h�r�憌�$P6��@3��&ؚ�6�٤`��0�q�fJ���JW�Pl�D�?�Kܮ	��j{p��(�|�ۨG�ٹ��3���$�xՎ�زI�Fn��=,i)�����96�xu��}~��ɾ��$�azt
���6�1\M��I�ڣ��r#k$ԛ����M�7L�B9瘮[�Y�VȊ������;Ϥ�beZ��e���I��Ly�#�D3E�m ��˶�����Xa�"��P^�M��=5�n=�Q?�RQ{�ޥ�w�"���E	LmӕV1��|MGb.�|	v;.�ꝝ#����F]k�?��ܕ��MI�J�M]h/Ҩ����5�C����!�}�%H,�-$�ى�Y��]�L.c ķ�-�1>���x�����J��XU[����D~D	���+�=��V�5�����Š�z�O�[���5A��p�I_��%�n~dl����֊|���=�����Qa�)�$��$��y�۪��ꙑ[}�����R,`/\��U�qBzl�����2�G��/U��y���[C(��c"r�[κH_�<��}Z,G1@l������)Z@T]9Y���QAٺ'�A-�9#��q��\��+�7�}�^Ӽj�+�J񁎤��6���i��0�a���o�qSK�m����:@�q4d�0��|��i]2�ML�� ]F����^�/�J`U���!�Ø� ���Y�,����uj˯�!�?"
;'鶞��܅e��0�9�Ò|l��ڜc^'>�W#�=��>>k��C���2����Z7ԁm{τ�%cۆ)Iy?k�����iZ_�u����̟%mv������lc�����b�X
MG�*``��:f�ǽ�K85��S/��Y%�ؒ-�ÿ�w���A�v"�3�7��@��p��U�O}��×irP�݇����[V	�K�4�]0@3Ͽ�1���I>b}���4���Y�#/"��r�s[�������XK�	� {~ߣ.�D�e�Pd�4�`ɋIO���* ������䞐$�D�I���L���'e�~���h�.��U�.���%0H��T�RQ����12���i�!����a�k-K��#��4�m�(:��ʒ��16��K`pJ�H����z�V ��s���ESܜ�`�?����׏Mo��Jk�t�<RT�LI��q�i����ZqO[e�ؒ������=�n���b<���..�[�E/����x��/�����_x+�*�F��"Cf�.��%y-���=x��˩6=&��(�T�5�-��N�v��q�_EO�*�T�\�E�Tؗ@v�"m ����k4SF;)����)'��Տ�O��=�%��w�ZU��#�#�g��D�������10�49u5b��:r�b�bYS�B�xȏ���u�rs����	0)9�%���Z�ɭ(�K]��I�8O<�\'��>�C��u���E�Y�����.=� �*G�!	\s�i<��Oݢ����ʦ^��H�U%�^m��tZ\�n.��t�Ф����\��AH�B���t���răq�ح,0�G&B�ޚ�Oi-��~���8?����0q�����3蟡jbql�"��T��'	�b�ǖ��#
�8��mo�k��ǟ��
ࡄ�I�_օ�E�Y0a x��X#���ً�?�*A����n��Ӹ��0��/��� �rײ��p���A��`B��G3>���0�ܼ��}x���tw��:�V����BC�4�#��C3�1YD�R��8%���(�w&���o�3��`x���泀�z!爃'Ru"���k���|���))
��Ϭ�qH�B�FjJ,KK0 em���]��j��M��ؾ�ւ�#��=�d��xEE�+�\J�5��%�+/��df?�L^�c�����
���.� yyF���եg4�+������;�Z˴Ϳ���X��La�=����z6�n�q���.Ȼg8hBP��C���(3YRz��
n��e;妍	���W�]�V�[�)��2��� ����L7���J��8�1�z��nJ�k�͹���C>���W���B���'���kz{g!J%��'/G����
2Y-��)m犸[�]���qժr�j6tS���+�p��UlT�nN���� h�&�h�B�^8�õ����R�@&�έU��>�0 ��o�m�Ũ�cM�DFBW��(�-�.��{\�$6���(wr��TH�5�~q��B��+K��X�
o�� �K�-�+w=�xh��9q>�� ��?Gbu|ƔR ���v�<��_vS�(��x4����PA1RT��� ��R�P�]$P���ǣ���o;O���e�9�{�-�<�W�fucd��8��d�dxW���3*Tk�g^ex@j1X���<T� d��k�x�ِsP퐙g�s=�فLZ5�X����3Z�s����	�[��=����9�\U�h�s��lur�(��e��s�&6y�&��D2��/4�����#��OV��������7�T��{�ӼkES��0�@q� �X�p����h.�%�г\I.�ު������9]8�){c$!oh�=OqP2<|�,��H����f �D���M����3�(��