XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��U����yGN�=s!�Qp��܈m��H�z6g?OTw�+#ؐ�~@��brO�U��Tf�\1��i#����H�?��"��+ Dߣ^�tJL�L{lڦh��ڔ8���p?��,�����v��Tq���6��^�'��K샠3�i@��t�z�>Ǥg�����c�q侧(ݭ�)��G��F"Փ:�%�&�W7n�s��4��%ER��a�Y%w�~'�Yӎ.�*G�:Mf-l�����H��{l��O�m,��]�$9���6睁�='����-L����n�Vc�@+>�����wm��Z[�腸�E�$�5`��+Ԩ�;6[�P����iG���h��Һ�����dx�^3)��|iTw2�G�'(ۧ�0
k�h6�hP��(��x���Xe�:���n��;�jK[��\����N)��f��%���2� ��3�Gb�Z;��z���a�� �#�!}�}��x����RjS��Q����Z��2��z)w���3��,�U3v�hB�PK���Ts>�'��jzjvڌ�1��Y��Zb&}�q|�_�5:��Dw� ��C�&���uK���OR�L����N�R�ʍ{�:��!�+�GԠ�>A��=4veE�uݮo� P,�-������N$���%��v�q��Ah�C�y�@7��˘*A����-�&�D�P�mi�b�iq��~��4��-g�qY�0EaTF5�:z�6߽�J��d�wW`XlxVHYEB    5e46    1530�����x��0���S��7[�tL?�$��ȡ]_��KP�v����DQ˜K'rX�yWK�I)U�:�-Tp/W�޻��;'hb�u��~�;R�}��:�n�����ߥ��<�Jѻ�Ƕ�P����n��iɵW���'��4r��Av:F�\�]o@_�iZ7Cx�~z������$��a�Bg�P%ٍL�S�Qk���r�yT*�"�X���<�MH	XV�C+ (.oW9��gY~�v��Će��Oy�t:�f�'Ґ�Wb�e�5c9<.a���Ƭ�+m�>Z������'W��q�P��	���� q}ch���C'�h� �@���2~$g���*�=�f2�RD�*tj	�?��fI!��=Q���8�4H�ܬ ~�>b��H�|_*�0=ⰻ��ڬ �������oL:h��\��{���4���s\�w[��#���q��^�HC5�J��"�b�=�ċ�o���a�DK�k�_�sZ�!����!�*}���ϫ>MUW[�@�NL�y{��;2=�M.%�a�NojS�T�߾s�kZ��P,�=�AR�8cJ6ew�&������߁�99�}^�^�0[sr��|z	.tS�l����A��_�Di�n7c(�"r$O�y���o�_�iC�)���nQ}�?w*0�^�Yq�����7�y���4iƲ�$��p ֶBj�[�B�U!��"�E2��`��Tla���Vh��Π�������gkN���a��E�ó�b�A�Ie�q32E��/��Fdyoj��G��q�%om8z���l�)�0ܜH��q1�Q���c��F�/����H�ƒ�";���L���;-����%x 0�7�4l/����;���w�G�D{�F�d��z!'t����F{ �(!0���3N΢��$l0��v���μ5&�;Ȓ�/FbK��W砅��ڄ��]s�n���kW(�����A�o�ؔ�yn�6J�&�#.��u�xh_�X�O�5A�C�g��+S�����t�+>#&r�7%���݁Jn��;�T<����0���u�'#���@5��\��̾�l�P��y��.���|GC��ivrg	� P�J��3F��3�Ɉ��?;����Ī�L~�	
sQ����3�a�w�^����ާkgY��z����e���zm��j�*�T��5ݖ�cr�Lh4_P?��;�Ŷ�x��R7��<{����k��[���2�B�gZ����-��`�wz�(��>��Q�<�"�������	p��xx�_ >�oI�����;߳k@.�U�Fx�y����7�-.[�8^\�y�~��j���xn�*�Ӽ��������RO�QK�+3T�Ẳ�%B�}GwY�:���ť���~�=1[K����J�ֶ��'X8@��_��h��Ӊ���cϑd���e�`;��RFgU��%Y�w�d����E�G-�?��DQ	Њ��#߮JƪU�*!�������A:�}s+�����y���LƱ�D3�ycn5)C��Ҥ�܋�蹈~�ː UW:��C^d��r5(����>]��%t׎ۚ���-΍�q�]�]�B�/��;UƠ�J���0��i��A5i�濸ɳd���#<5E3�j�[�Ǽ��Z=��m�j0�Y7��1�C"3�J�5�� ��Y��wN���si�l$_�c\H��"�4eǞ��xB�����l|���5��������[ )B���������mo�Ԉ%9i3��՚q )�D<�_0��D۵�$[h���"7*N�K�F��=Ɠ(|��D�|�T)��TE��L>	�.�p��V�����j��t���#�7���J�y*��	�1�K��5�c2�T��k���c�C,�m�O�T���߅�B�V(W�E��8Q�VG�+�uy7��= GUϢ��F��ЖW��\)������M+aF2E�]7=XC\^�!���
����u������Z1�{�I��JS'4H�����ئB�sLV����\�kd�}�{�On+^q�ߕ�X�UI�<$^��,��V������$V��~?���C�P%�h6�Uހ:I�`?����n���)4��d2߫O�bY2�i���[�iu}ǳO�vd^6R�����r��W*�|(ր)'��Ϫ�}��+k��`З5y��"��^��K�PDő!�/�j�!�E�|�����.�T!��OJ�g�����ݫ�6��+I���x�~�uԂi
<Ն>X'�iG���8E�N�Tu��2�X{?t������fVd�V��򗒳!��z���
��߼rÂ}.F�&O�N�d��Y備��3��k{��b��f�<���z��d������t�/݈�&�H%S�x0V�°�K��0㽠!c���� t�-9�Yib�~�D��tW�5>t��+.�(	��Y��hɶ;FLƏH���lm3B*�J�U�vy� ���ݢ�
�9`fV�0chrs.B��y�@�?�|J�[��'I���$�d���%���:*p��q@t��wn˴�V���R�^�O� �0�7\�8��^t�Y�3�*���5��_�wm�%89�yJt䠊����Z my��4���
�� L�F��h������}�����0~?��5����0����!a[@�ڊ6ۆf7kL>m����lU����ի��a�V��R��@��:Åo���/�J1�a����ggB50/���nH���,�B�:�J5��������t��fq�T�1�-��o���M���o�HԍTu{�BQo�&έ����b&{�;��*�5�ڢ|��-� +w �[`qઃ�߽�@���R;L����"��Z��@G'x�>�E���e�}��"�zwt*�[��,�]��Ŀ���l�6��V(��{�(}d!h�b�E �뗡��Ѡ&�ɥ�dw���i��H�Rf�c��p�)|��o���ѩ�3g�l\�i��q������=�eyG�KY�x���N�M[Y]�����p@Q�5b�3��7�Y�j�w1.��q�*h#L��5;���ܟ���F�C��,�5'�%
�����7?]����/˾��FCP�C��|}���z4s�!^^���(�Q|+����a��$���kC�-�<������&�/��W���ŐӪ�W�����^�����Zq��h�FԵ{�b"ߑ8�d |y��R<#��7�?�	���ڔtH����`�c��c�A�&�����,Jx�:d�=p�|IfV\���K�e#��m�Al0�)��ZcW��>�k������+�������/�4���;y�����3�~�[��p��s��mm�GH���6��$) ��K�� Q�_�9�A��~�8�\j�/�3��d�.��ϙ�Xc�E��]�|2.�����@�v���6)J8=�m ���s���tY&��Ԕ���@�9�S���֓���n�}��
�ƀ�[������^�t:TN͢˱aY��C���<8���vTL�É�A�GcY�#�6��Qx3�3��z'����E�V���9�c��~��}l�}#;�)sfk���i�()�	j�ޜ�m�g�A���lM�؇~���K
�j
�u�{O����"�P�	�?�C����"J�+��\��8��H�ʜ9r{�L{�ᒣG
�|�
����=�Z�����]�#�a-Χ �AA����>�ǜ����	��i�C]�=�)��Pr=4f�����d��e�C��[�	ߕݻq� �5N�-�Qq^��G+�F//�0�ϧ��O�vM���x޽$j�Bt�<�l�=x���c�';w-��hp�
�{�3d�1���!Ӛ�BA�����4�ȭ˵���"���⁁N���&�ۄ_��(����-�]"�~S�G��`�+a$�X��Hb�E{Դ�#"�ȹ(,�������͏O��������2�
b�~�=i�_T��w��s36cr�#���ß�!D<!�F<.|c@�ko3����9�&�<5����n�+����W_��5]�
浿�����N��ʨ峀)���ǳ���1o�]v������Z3{lm -+�C��P�܇ڱ���6���7�� K��E��k����#�*(e�v�����/��s� ����f����X�_���Ģ��Vg�d�ٓ�ֻ����HA͂�)�j�S5����?�-~�i��G�11�\S@U��Ϻj�_�P���ŷD!�*��J���a�O`��6
[�,E+�D;�4�u�=iFl�_]����q鶸�gl̓���T��1�+
���%�-�,�[M����T����@6�Ӱc�t�r(�ܑ�N� Ym�Y��Rc=#��5�;�S�7ro�Z�p�=s������4��������_�c�A ȰUfMde�WK�,��P	�ݵ�/��I�`z`��y�����-"F���,�w�7Q�d�F�ر���ll��ye��謻��i���jIT�+?�v|ś�ڠP���m�M�hGt��+h�7t�=���d ɳ�����}`=B�n�<y�����zk־o��uL�f�v���K�����Z��)G��c�������i�M-ܫ7�G9(�T>�#G0!p+�gc��
�����sk�f�������v掮y%n�K� ^�0���`���;���i�wK����u�����p��.a����S��6kк=o�qR�-��R�ǅ��9{VZ'sLy�kb��,�b����\��vH��Z��/Iw�Ce��a�vR{,��қ����!��y���ЩMr~V�*����\P�[����;s��Sג1�Pl�rOi�����C�����Bt���k����G�Gq��[{��!S�]���ӕ���9d�xm�1���G��S�u�]e��Y$������KC�𩭣h�P��[�^vuG�J��לD�x�����c	�s��ۊR�����d��Y��˖+��T�s�"tyfk��lg�������u�r��t�,��,{�g���������)0k�[]�e�J�8��.��w�=h�S�Ws�����C+~&��.�d7��C����k`y�݈�ذG�7�ϛnOx��|� K�k�n����.�����7���[߱Q���?ŧW$tH���)�l��¦<�Ϊ�-��+� :�/��_T1�t��	��?zQ%�F�!o�����CN������o$21��>���ó�!����4����\�Ź}���HMG��K�:m%^��1�P<W��#CS���c1��4���ȒײgF���璉�9�>�k��#Ĳל��=ͮI�16��^��� ��|3��� ��̖�\��;�m)ɪ�Q�