XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����y^��4�қQs�B'���7�+TKZ��G��;�.���X�U;r��bq��pR�|a0����§���rگ��LT�J#��Dpzf~t�.t~�P9���J��A�]K5�T�Y��K���m�+;
<�Cʬ���h@��D�(�Ԯ��y�PR��VD�����:�JR;��r!y��F[��2]�v�@깡���1,��h|�y�3����h)-�L�:���6��~ CT�t1)�G*b3yH����->X?��/��V�H��I)���*#k�vo�󈤾�]L�ڞV�������I���Ө�a
=bX�͕�Xq(T��˰̰�cHE��谭�ן�-W�Y����?�4�;��.��D%�� �Hإ�2�������xTr��Q�+i�Fj� �-�Eʩ>��W\[(�Oɛ1)����jr��K�χ�ox�?��'[l�/�X�׋����p;J�NR��ɠ��r����N�v�	���q�b�i�u��|���l?�N춯�nA}h��S�dOs~P�_�m/w�V�0�wk��O�3*8�����5��d�Af3��[k�$�k��r��3�i�뎓gj)R���g��K�G�!�jn-��N��ȁm��|eCɸ����+{ךԀ*v���t�vt�QQ�y��|7���~n;И�����8 ��R��
0=�����4ygG6ّ��՟'r��}!��ъB�0�����s������?7���'bj��(�gr��ݳs'VvN.XlxVHYEB    fa00    2910����k�Z���pc����!����2|�쫷�p@#�6��u+pA�JJ}>{�֊U�^O��Xڣ�~i�˴?��L��i�ǉ{e��7b�~?i*_�A���!}�&�z�j&�S�2�eODX#E�5d��nR�ʔO�1iNqF)��;���>ө�������|~[c�2bn$�[3����I��0��p��m
��9:�|�ʇ+X�]��C�<���̩@
�,�,"%x�{�S�$��:>ЌG̈́�����DS5գO4�v�ZQ���ڝ�T��5�{��\�\La�sbg/vmS��k���}\@V��EN�S*B<?3���h�_�@�ur����ݴ���l���k��Ǯ�2��}0�_�_�Z2�T@�κ���Y:,?Ә�e��in-�=����7���r��9�R7���6�Ǐ���,E	��C��2,�Nv�U6h���\�9f��� |�&���+7Y7D��I茞�E���IWm���I��HH]Zj��a�tR� ��77X&�:|�q7��y0���I>�`�tq�.bJ��1��.���UQ8^��i��q��a�J�)*3>`�UY_�U��/�1���e��Ԙ:��af�c�|/��Ŕ�B?S��$6z�([ �~o/��z:��}��+�	,�J��2|��y�U���������4t�WIa֘��d[��Yl�ymU�@.�=�=èj0E�v�|bM�Al�2��<Ђ�B�(~%c��=�(�4��T���	���1g6j��B��b7X���T�tW�8I@P�k��%w��V!6^���<�&��G2|���0�J�3%��w�=�5ե�p(�����I���r��[�*W��.va�M���aR+�Z����"��͡��L�W6b�=��%�u���O��j�L���^���9Zb��G��n!	BX�M��p���xk���O�<l����JixX��5�^Z��O��ğ�H�̠}���VᒔlM��<��0".�'ʋ�v�?�%�u���9y��M5I)��Q�n��Ȁ�N���!)
uQ	v���~�4�Dϼ�ra8`F��U$�"ӱO�u�{�����.����1�� `��J���]m�����t�A���t�e���0h���H~~	%��[([�N�r*&���Q�h���;�o���j���SB\d4z(���:>%��Z5Nw�*�W(�N!O6Ec_�mڧ)��>��4Rgrۑ�C�a�HDQ;�1��=U�?����
�j;�R<R�	?�9l��'۞W=��p�� |��1;�b;�R���Ml��nD̰�FP� ��Y�~	�;O,t;jp�u;�wa�m~��N���HR#̾P��2S%�,�[3���,��ڰ�xD�@_C
���j���e#�L��Ķ��k�ɮ:���<�\㖲�Q��*F���~̜\T��r��K�e�^���~T�`#ʞ��,��Օ@3Dа����6���R����{e�gx�(���GL��e��Ih��:��E�+��Q��kH5�6�)7��s���;����@�.�ϱK:b.��|35&���p9�]�ܝ0���w�������[k��:g�O;VH:8,�f��hPͶ����Թ'�gE�՞�W�WQ��-D��W`�y��G��J3��a���(�-�F�;
��:�1���%#^l��:��!�
�^:��������'�b�#������q0�?�uA�c����Ռ��b�6��Kt�ꑺ��L��R�\��$�S4gg6��X,{�є(�@+����=.<J�zG�����s0����qD|g��M~?�>�I�"�l~�~�m���\t��!�&ے�F>Ҏ3^ձ���Er�ы�:�S�p�m��yD�X�{a�,,� a�P+��:f�S�|g�?AS�o��2r{:�����1u�y�hGb��Q�-饹�{��q?!z��Cw�Я0�2��w ���=�b��Ϧ������].}�c�He��L4���dcL�\�'2\w�v������;��?M�ћ������С����:<�ж�8��z�k�T�����W�5�6�C�����	���Qp�To�lT���H��I�c�����1�u7>AK�6�b/O��y�����uB"�����sS8���t��u2R���`M(��7j�N}��Nj^�X@B���-��ꁿ��ukN��֤�>�Y����P��g����~�XV�a5������)��׫ܘ68J�5_#7��e�ɶU�4��9���R����4�Ex�i��e�Q��1c9�b���[�4UjQ���W����n��!�%�y�<]��,�8��)�YΔ�p�7�x�y�X����.�0{s[�V,����`~�+����b9�9�x��T@�㗥u�OS�OEUuˎ�g����*\������-��q\	+����R�"���fN#TN#bM�W���\����:X�x��Jn2��:6�l�-��
>��Q k�	Q]Ҷn�.� �c$���7e��$�OI�BJ��F� :�6���G�Z'dťEG�+�����Q�̔�(�)�J-RO����#ԟ�3�c�%���@eo>�>��4�(}�U����xPNd��&��%�D�Cd�����y���Uƚ������Im��Z&ѠhP���'5����?S8��5�g.�`Z�)���9�`�^�2��ԙB�)��%�3!_Tc�.���@z��s�c�!���b=��`�EH6,�v"��_ET���������Pg#�[��<�ٜ��3�Z��9�%')�U��8ä�&��g����(��B�"��CL� �[$�|ά���7��*e�[��/jjN-?��������iS�@��P��SW��
Q�'�.8���Ab�q�1��p��Z���;�M��tB
�DU��4$e�]�F��[��'K���\�E��4u]0p:���rm����6H�* �}���Yۃ"���O8��"M���y�+�ƫ��V�u�a�{R�hX�	o�)�n�>[�|�J�b� �rFnD��8Y��^,߇X�፱4fo��!]��y�5��I������d��%���/�w�<��6gX�� ���r0�T��ƀƇ�H�(���5����gQ��eAb*7�&�8P䮑���j�j����p����P�.L5U�H]��TWezإ�$�v\���&K��i����>O�FLpcn12	�M�u^&��`�N͵x�'�����:F�2b�F7O�̢��:)��d�XI�~2fIK�'�K'���wJ�F�X��
W:�5N�2M��Q8Y	����O�"�_ԒMa��Mʊ�I�Ϡ� ߏ�Ad�*IRV ��g��.��-n�l��	�8qs�Tb qŗ+-|� X�*��X�y�,���f4���S*�%�ݒx��v'N��p9�*�=�a�ZIԟz� �¾:K:}��ю���u��V�x�ʗ/ЯE�]��'�F�͢ԕ�ofm�n���1,��v���ʳ�A&љ�a���ӞZ�y�}���Ӥ
���(e~l��1>��Vo���Q��n�%~�89�_Gq�5=4�W����,b<6��;���i�P��z�˛"���㑅IW�=����E�q[��#H��7��;O�y��G9!z��hF��\u_,dȵ�}�CF:KD�L��>1ߒ9|UKc�;��8��֠Fh��"�@�$Γ^�T����
�f��߽^B��9��&���s�q(�K_�a�e�Z��W�5 Խ�4~�ox��*I,9� 4��3�֫�y����f�ο�s+ ��D>MLȐ��<*�4 :��Y���Bi��-܁�,��Z�"h~t��qg`D�`Z��9h�W�b�e8�.�	Hu+
`��參���9"���^^Ԣ��N`ю����y��s2�_爤b�qv[�C9�{�|����*h�H�t����T�$D��`9�C�V[>���iw��w:��;�׋�Q��8L5�I>tLR�c�\��%�T�XC8��(5Q�śMR���y&qJBa�ԓŤy�9'.!2�8�����.�D�=o�I��],I�����i}�^���̗�q�Q��~@��mw㫵%���H�v$ZϪw��:�5<޶s_k�8�m�N1�����[���ߋá2�q}.�����^&Ry7��[C��'f�\1B%�\�r	U���|0��Q���,L�m���/'|}�¶���1x^�X�e� ��tR-h컖
��mK`�eX��2�I	c�q�]|@�?Ȱم%�v�E�����,����x4/�_��T'�ĭ��C����+f�p�,b*.⭏�H�0��S3��rY\]�j�Il�*�B@�R�>ց�������.�l����Pc�֖+�������W��vz��͎�Bg�2k��p�5�o�םi�=2�g=��vPm"Eî�k�MR�h�h��+������<lJ��6��wv�փ�����C�-��ch� ��3�Њ�2�f����@���D[�e�Z"i�`��l��{�!���kO�|��u_���1>�ӧ��^�x�%>�P�XD�BcH��ך�X�K�.�YY���b��8���Q���r=N���-�ȼ�掲4H���z�\!Y�`VH��i�>�t�Ѡ��$��g{8�Ԫ$����z� Lؿ�LF�����MPO�>�܌�x�U��c5,�K��~�<��-�e~���łfGY�m�b2/3����S�<����X ����SDk��$�ޙ��%�T
<*��я =�T�g-�:
��5�_nt1F	�b���O��J��X2԰��,,,��'Z�6���Pcс�,�Sz����l�o��:�&��xtJ�{Ȯ���׽:����=�#�Vh��ߛ���ݜ%e |��Ú������\��ւ�{lZ�-� �9��m֡{��) ��=�oabF���{��k�ԇS-��*�~D���?����l ��Y�?WNS�Rj�"z����D��r�ާ� �f���ȞW���,Ձ�p'w�v���O�:���?;�tѹ� ��c�}��"p���xf����ǟ�C&�e�e�*=����	)LR۸"ݬ�mM��z� ܵ��jGR�~����$TFa�@�YW�B��{?�����*	X�s(��_����4~�ן���$����.+��׷� 
�`G�ϡn�=�f(�F�gqAJ�3�4��yT��8�އ%����ye���[�	*�h�>-��:G?�2�� /�,Mj�6����c'��OZ�:�5��T�Qa=�&$�h�=��Y�.+?�)�]������! ����S��5�?��w͕<*m��{���4W��Q�������=M����D$H�s�HIWFA*G��3�8���fs�=r��im���]�i�+?��_~N�!�u�j��D&W ��9"�l��S7]�c�I	q9d�Ug;�يSSB[%K�j��{oڒs5��������5̸6D����
Z6�5��@�DXҺ��|y��cn�ߴ��~��p��*��e@X�eNX_�]K�8e���L~-�8-z������jG`c��O̅�3��f�rSJ�	�l~ft��mBG�{�+bv��i����9d�\�w��qs�
8��>i���'���cm����(h`,��"^־��<ZV����rH]��%�wQVK��;xC�DZ�aWM����'�~7c�T��+��t��ki�ld���s� �.=������0Z��5��ۿY�b
[X\�gQ��!.5��s2N$�S�h�#�i�+`	��'��2�]������a�A
�`s#���s�ŋ��X�$�� K71madڍ</q�WyD��w9TFu^j&!�׺��
<��=D���[�d��J�n���`���V�c�#T�T�[�>BF���N��GX6:��Ʉ@���m淮��Y�W�k�S��h;���������ay^9�^\P^��B9X���7�f�Ǐ��u�z�)��X���g�'V��l����,���j����D+h��1��g�7�К4�	g����)�s\jY4���j��O�q7��;o�nZ:�4����:�`w��08��|6}v�ܻ
6O؈��Z��U��i� l�G�r�1 )j&��%�*�l�1�S�����~j�L�~@�x]�4%��|R�oUe�q3����@��n�_yiEu�L[9����Y�Q��1^��p��.��h������wҼ�"�U>�<�~���rM\�-Ċ("e�6���?9�ݮ(= ��?�/DИ�Hպ�-eJF|��as�(��_'��ڥ.06�[�&�Jqc�L��]�!�N�Zj#/�a^7��!���m���G���{��R����2x�(
�ϙ��|�Ö�`3��̇�P?*N�/-�����*�9���!��U�/�+�(�&�0�]V�*�!���e��iOª�ZE-�Fx_���{���>(i�/>Ƃ^�V��9VxavJ��`~F
�66��':�Y�=$:$�2��<&%kB�a�/���<�rd��-Ʈp�*iU��ھ��XEZe�^�kB��8~���%b\��������U5λ4���������2�ձ���)�ã�.XS��g�b������^��:B�ϣ*�,�?�������׏�8<g�5�mّT�	�=t������\S�z�,��h�>� ��t$��2u�j��j�����x���v�vH��^t]�z��ӹ�7��~^��|���if���׃�6���l-�\�4�i����g��(Pw�͑�
T�����,|�rɸ'Y3nXP�J*��${xY�-���_�0e�5K�\�V��=ҁ�~djyŬ?�ZE�"K� _+��Y���1�]���ߏ��HBZe6�H�6�yX[��u�?=��ʅ�}�u�c�5L��� P��梼�E�k���GH�>���yݜ��tB�lcU���ڕ-R�`��\�=�m�3�ˡ�	�i'�Y�	��՞�Hp�jAB�C���ܙQ���)0#]i�Ty������	�}}>�CLN���ub�$�0�',$'��!W�� 0�v��Q�i2�a=r�jhGl5��Ts3�؁g�9���ٿ��� F�C:�!� `]����@�"vX7i���������(Z���������z�T�g���&B�x�S��_v$�ɭpN�'�4�ˇKs�h�!f�>���;�?���0]w+;��.�#�|P��(t������Lכ;����T,����.�se5�rQ���tpF��9sBV��I)���x�#��|��ܥ�ꈗ6����}~A�ͥBB꼛;6
�Z}�h����i�F=���W����%e��cI�/�A[�����-f=ؕάj��'��nZ94�?������P���9��V�nlrL�z������!��_��+���Z�\�O��=��yø�o r��d�sb,Y�mdi#j�ϛIfO�HW̬����S� Z�E��;:��S�*h�Q!�0C��9 G�%��7bۜ*ӊ����$�����!�g?�'7����8R�߀��_I���Z���4q;��ri��U�oa&9��r�I�ZYssK�����9)N5�"��;V�Z�A�[�S2��O|�n��jV�p{�ӏ�l�?�pIv�ϵ/���\�g�QToDT���;�H7�R���~�g���Th�"*�lt��,�r�\�il���#��j���}�ɍ�k�?{�C����������5�6�.%���c�s_�U���do��F���F��P��2g%�dX���N�}�h�s\��8\C�x���$�~���]�a�m���m���ۘ��[������؄M������-��ŵCКoF�碫�kU
����3�x�0t8�6`��0�T?��Km(@�F�*��������0�T����g������";v�"��O�0r���`��� ��qXD�(!�:��G�9.��iN%�3�l�s�+g�t�?�(l�VLyb��le�
�$����o�v� �Q��d��/#{+ܡX-���pJ�R�U	&�}���Q[>rV@���4�C@Q�ФJ�8�Gz����#R�u�x�{ur-�E��O��?����}xK&�<jڜe�]�(���@�eOB���Ìm�G�oN\&v�
$L,}6�?��#M��� ��z��q8!�I΂t�͙�z�<�:Gf�h��_f�MPb.-�{�v�>0�u�>!W{`��@y��"���ː2��x�_u==��F|�gL1�:�O��)��~�$r�zM]H��ʢM���s��� �"8z��8 l+��s��T��F4�'����p%�d/t�";Q�g���~����Jʂ��p�ES�a>����_a���Z�t�;lA���@�(9F�����w�ixI�~�:��\F�~�՞��-sO�5E��=�)��)�H9U���V�f��^8x�v���k[�Mg:�x��ʣtx�]ͮ�"��{NT��Jܞ���F̀��*a%��Usݘ��Z�O��>�uڂ�m������o,�K�r�p`$��!SI������4�Ԏ�1 �~�T͌���M�E8g�v��w��5��F#«�Ou�ErV:5K%I���ı[U��o�=8p��xS�s5�1	�����a}c*6���%d�ݟa��P��	9�D�q�z�����%ާm���	�([.�^����p�
�@�/��M�APۜ�h���rW��/l��yJ%�;��x�ye��U*�b�W.@�H#�������,�� ����Q{#�gk�ѭ���}�*���4h@���o"^�N��5T����O}v7<�v2��ج�ׇQ�e.���jG�,G��0�ri�Mɥ�q�p���d=�ʏ����k�'@�Ut���^u|?�'Q�s5���߹��|0��c�s��Q]�G�F�!U�=�D�OKsE��Ӎw��~	,m��W����dk �ǙpH�(Ƚ���lf��"���TDXZ4�����u��,k� $m�Jz����%��R�@}��v��3L�M��绑�(�ڨ/�K�5�8��x}����x
�m�v�&<�����ݺ<6�[|Fzc�+�B�d0���+��:O)�ޥT�6+BV�,ǉaG$a��`7�E�~!y���'�O��z���n�g@���P�L���Y��sx	𓕕�Y���0	��27O�/Ȼ����Fq���r{��C�_�������U��	#��cU���+�D瓇��
�Obm����`3��)T�=.b�>�k'
N�F�-�$�"N��R�K��̩�&-5<'r×4�Ş8^�bB�v��Kst����F�h����c�$����\{������)g�A�P\d�~?�e�@4���͹�F�A����y~�C�-��p����+�ѕ'�3K��r���1�'��v�vV��0����c`��f�W�=l=i��S$�#��t�3���z�|c�V3��{���,���V��	Y��4�M)q0�x�kM�lQ�����x>�xW�ZP�p����
�8�{�4H_Hx�0m�7��K:fSE[[ߖ�\.��Nj �d.4����8O���%��t؜,H�S0�^rV�'<�ςّ��*����a���W)�~��k1�x#�2�%O�� 6%�J4
�b�%�PnI�"���xѓ��6�պEp��� ���1RCn� ��5�V�H-NB38�MD�!_[ί����CKatj�����Wi���
d	u�����;p�����򔎋�H�d��&�Iۃ�8(��mn@yp�&[��1+<���}���}�>�ؾU���C�1E��@^���5h�Y���T>q%��k]�w�DN͘{��� �+7$�Y����l����4q���Kr_8���%0�4'��_vi0y�x�d? cD�=�k3���$	|�d���Ŧp0|�]�N*��F�n��!�o@	w�&	,��M:�_&��f�����9}�='z�Ηug�#�3*O���RPsJg7��j�py����v\� -���V��ݜ����썺���.shjs��\Q�î��*��D���(�=�I�H�S�F��$��0O)дܸ���']< %�`!�R>�B~f��9'oVXA]�<��i�S��L���bn2I/�&+�!�O��I�X��n��� Xh��?���cZ�����-���,��y��]��p��4�-��,e�Τ���/)p��,|R�����R��r�M�]�$6�ɜW��x��ʊ>EMD�Yf���w�G�Ф,ܐ�?݊�����x���x�Y$dՃS���vXlxVHYEB    6184     f80F�ҵa�j�5C�d%�3
�k)AlƮ�a?��i0;D��űM�SL=dT �_mʢ���X�\�;c�[)
�_����A)���Q�ܲ�]R@B�i�Vb�T��ѥ/b�sc9�
�5:��w�~��ѝ�)���x�&��Kǘ{�}{	��[�_] ����V �L�rhKʖٞ$.��1�e̎W�I*���� k��+PM��� z�_s<LG���K%��7�����I��`q����vr�4f�]B<��}�'��nTq?����G gJ����3k\�]K[Q쫱8G�/���!�����yE{���Gs2:�D��#1��p��b!��Ӻ��2;��X{e<M��G�(�CѾ��.�l�����W$n؜2��4�ɑ�#� �,������0�aR��4)K��g��J������0��m��)�Y$�K��B���2�u�0;�itW���g�rج��\����s�
h| �*5�3S�%ˁ��2��.A�n����Y���ʎ��8`T#��G��C�G�6���ʠ���Ǒ�,��+��W	����8����t��ɽ�R�	{qߠ=ʭ���P��R�](V����w	���]
�9��*�C�d>�����j)Ĥ=S�BM��6�(֋RC��q|-ܼR$�D܁I��4ݼV��H�ͬa��z
0[{��g��� jc"����QǖZ�*�G{�]�3�W��/  ~�F���z�+�	Tڡ��lc�܏sH*����0���pD� ��Px:��WZ��rz�e�.�o[��i�}��nr����Iv�+_�p���~fN,o6U�I�����=�$�jq$N_�:�Z�"��CO	�|���c��1-���CY!��$;���7̐BR�~xl�@�3' �bE�:Td��_ս#��[�/�0[w���d�&�]RD/�6~j�xY�
Z�^Yt �q�'s#$�o�If���t���sL��$�~d{�]Tn��U*an��3�LKt�.�jϐ���TE��~�C.�ڗ-���WL)rz!v-}�U���㟥U`�E�����뚗�&��z"���e�� �+!�?N�x}l��iǜt�HNu`���ގ�9�����Y	��b�T�C���ޛ��q�\��ܼ�"@��ĭb\��R�5���#�G|z�^�_�����@�u�����m�6�#��,��hP������F?������"EpZ���Gڋ�ۀ;nZA4���p�h�!E�р�wږ�2�ka�\�B�B��ݎ7���^ˣ"T�QZ�ڠ�|i5=8�tԎY2c4-�^�&^���F?Ae��8�y���D�Έ�ȢÞ���������:�o�0���=Z���A�H�w�ot��w-fC!�N������_�-���p��,�'��|���.����;���k�dC�;.g/���J��m��3n�U�E{{VN63� �Ǥ7��l3,�B��装�4/�>�+ԍ�I;gzᚺ�=�[��ָ�&9!@�<P�����=�t;��X�R$'pY�	�V��6[���:+�S򋣈���y��˴�+����^L���� ��PʑVH/���N ���W�/�O\?���;I�q��nN6S�}��Yܟ"OV�L�oVM��s�
�;6J�z��GX���u�+n/����K���ǻ�it7�yt����y�7���&o>���;~�O���
P����s)��g��ϒ���Ѧ�dnsp�P��W��G�l�gW8:�́�]l�`P9 ��|����<�7~�{��â"C��q�Q8��J�ÁT�t2>��w/����4�N����_��3�1��.�5��K����2�w0�-�/A����׻T[Cv^�Y_ך�	)���c��3��>5�e�\�"��+A��
�1$0��;��ytL%���J�\Y���0)ߞL)֙]3q���6����v09�m�B���X*\/��I�b�!�1��h)��y�sb��!W������H��,��ڕut^X��-h��w6�[����CV���/-,��_
��P�^_��)��#u����(�r�b�˗평A#�u6ZhL��"XW�Z8��ؑ����չ���SUun�a��Ba�D�q�����4J9��u�v�(hc�_x��E��<��m}	��@��A6��.3�O�`?K�=��*�~��,(��U�{P�m���C�!�t��ra���@�[R�b�����Ej��0Gd����� �����-i��jYF���A�at�?	3����{����zh+>�J_�%��}�LM���DTd6�6I�x�y����9��qs'�O�jÐ����@2ykPO��k�/��r�Ǎ���!�XmMǘ��s�2��Z�MX�֐8g����5�����yG�MGO��i���S؝���!m(;�x�Y0ܵh�:5�;�\,[�8��t��Y���*O���Z�n4ɏ�h���~�O�� ��@�����'k�0R �4�;4�=EBN#T���Adp3&���9N�.�/.���phIy�qVд1���<���=���ú���	UQ�>�< ���+�W��������id�J���P�*�zOk���'pr�m�f��P"�@C[�i�.%�&�@y������7r�EXg��<�]<�b�j�K<T5�|@*�Q�;���tŧ|�R��+�ǵ�Fsqtnm���y
�m�0H�	{�����*���O]��������H<�9�/���8���[�gJ�Bs��ya&��c��w��6�>at�/QnL����e�j�Љ�i�z��j�s�a^r�%��K� yH%��5f��B��=�!*�>CB�?j�肶Φg~��x@R�`q�wd*��H.]D�`��|������O|]�[,0�ŔFq��U4π�.d���[	���=j @��f,-�g��������A�mH!;*���M��M+��^-������4Ġ�DɜoP �N`�ެi�c�C������y.���V��JX�ju'�T&bA:v��_W�S���Y�*;f�Y:�R|�7@�?�fm�����xq1=���dӮ����;U;��z>�Ut��P�X-�ڄ���Ax:���������o[�I����4r� �J{� �?�!�\��; �@�z�)lq�_ٓ�,g�A�Z$\O��ڸ���I��_7�=��d&�l�-$c�
KK� ^0&�a��ۖ�Up�H��`�Q3�w�?��~���^�#���.s������i�{�A�0教�>���o�\Bc����C�?tp�d�������ٻ�R��r���9�O��8��ʺ�:�<�b��r����;�
��t]PA@��^�=ɴ�3.�l���c��J�1�T�/o��0�J���Mf�<|�����������\RD�.#����3&�OTs4 ʬ2M�L�3�<[em��A�4��`�Vk�1�w7����Ry�bׂrJ֚��lv�G�V�C3��H3��s��|�h3�z�*V�� �P�F��sem.]*'X�I������X>dR��L�����`���e���4$ʅ� �J�ݙ� �t\7mK���-�VG ���A�&wC����V@�y��x��R<X�5�������:�h�����=�d�~xp��d;"S*�k��k��Aw�1�},�vz�\���<;&n�ڙv��š���������Լ��;TD����.
�4������?*ρ3���2o�≢��;:�Q����28�榏�֨�}�>I@ɟ�0W�t�y�\������p<.	���OŸ�Mmi���{2��@Ϝh䛴����+���2�f�Ϛ����,��Y!z.�Eh�e)�[��h� p[���!~�h��+p��u�"