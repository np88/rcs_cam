XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���@ּs��{M��[�/kJ/�ob��ؒnH/@�Ji�qTVw�rP�ⵊA��j���f�;srL��P�p��[�"�M�{���-�1E����ȥ������ݐJ�̤P��(B	?R�� Gh�Bm��ST��xj�R� ��5Of��E�ώ�����/�+��崰����gU�3�T^�[���g�~��mS��å���hRw5�� "�ۼ�~�X��E��n�E>YC4�B.㐍YG"�z�m�N� /8,>��!�\B0>h8�_ҿ�fbH�5C^�$�F��+���)����O�@���20����S�}�I��2��ŷ���vH��ca]����tܳb����P��F��I;��κ��]���.����3N_�!f����Q-��>���|wF:��/P��Nsy]�.�o'[�3Z�=G��$9�xh|�Q8���#X�0I���e��7%�R~�ֽ��J�z��K�ڡ�v�La�w���ъ������K����[�8K�WX�=3�v��U��K�,L,%�N���L��J�WL�L �+���y�0��w�p�BXj���%�5�O��@��2s3[gG��'#Mb�;����
� �,��dF2�ii�����8�6?pz`{�|M�������u��I{SO�L̄6�%T�	q���q�ZꄳR���
�W=s#�ڌ�j6Ѐ��+o�Y���,�m�^�B�8k~�]n8�$�D*͵O��'>' Z�(	�c �*�-���pɠ
r�er���vXlxVHYEB    fa00    2910����
���69�֡Y�*�\�k#���O�H�\�?����փ�Ór��hx��P#P~Vi��. i���a��յ�	�9�K�D�eP����Zz;b�.���^o��v�h0����Oo�x��q��3;D}���U]�}�p讉#r�7����I�m�8s���V�ټw�ck��]��E@���[F%�d�W��Xz���'(�w�k �S��Si�{d���1�u$B@!5@,���O~I�_�����&7c��`�<���&; ��%�0#�%#r�/��/��x��4o�0sSY�%q�Ƕ�wwW���%��UD�� �v�Μ_�|˭�хp\N�f��»�&�si����$p^My����oi90���\O`��|��~�YH�#׺ v���d��$��]�yg<�U���Jmҽ~�%\T1�EC��6���8�� 6񬨡�|�awT�;�fVWA����#�qv�ѷ�M�$�.ɹ۫�L\�p�Ҍ����7Ƴ��!nt ����cf�1���OLcmVXJ�c�Ϣ�btB���6N���照�����=|N��ow}6>�_v^w�K�)��J`��e`Ny��ߨ����o�� ���j-B��{�b換�b��3o�����Ύ%?:�fq�5��!7	�"3_�U�M|�ƍXͳ8��ɭ�wn�to�(��֐x\����>O�=�j��v�^����)����_K����s�@�W��9�S�+	������|.4L>S\��C�3V8I�_���'��P?�lpX�bg����s9x�c����7%���EAyM�a$3cH�O�z��_G_Y�0��p#��n<e �����Nd4p�ccc�砜e�:s�Ç�>�����40��4l[p
��;��9�C��5v+?�7W�,�FF�3Ry���	1�ؙH�?�ʺ������L\a���޽%Q�s/��2����7��ڈ��M3�m�/�sM	��~�>y��{��!H'�U�7������j\?��!����x��ЅW���G��۠���C��ͧ��\9��Q1Zʁ��u�^aC�)�.�d�����f1'.�_�i��Rm��h	��n�>�K�G�+���P��}��v�$]��Ҝ � ��t�>�@^;KY�G�w_T���m�wT.�ҊC�z].��谽�F�.1����ƞ�NϱQnzx�)�(^�1}�H�Q�<�ir��%���䚍�7�6��:+����%��-�V��Ɖ����~�j��E�>����G?}O�$���-�s�}Kq�kg��ȏ
V<���%��f���gEa]�brU���&g�n�W�J��AW��ӌ�.-������(07��}��y�zzv"Lʙ�u��`a�#D����^����Gs���x�%4�^�X��C{�U �Oa�+L^ǨRpz������B���u�^��P៏�����%����Wa&A��W�\RPb�_ �nX�����4c��ڄ�B�xJAxr���X�sUA~��)�v���䚐��u�}�w/>����>�tZn��A N�}ۈw�c��9���%��呟a�B�!������r��H��QB�')�_8*�Q�9�>��E�.P����W��`'��^�e�f���	�h����H�(�ޗ��-�v`�%'Բ��b"�:�^�>Y]�6���Б8=�����E�v9�d�$�:>H�4�����Ttܳ�?w�v
�`U��P���VXr�)�p6�A�C�3���
���q�aZ������di���x�*��C"H�=z��NK���,�S�
o���Z�G����!v��:�hL�h���`J+\��M��Ѝ�}�����6}�;	��r�=՞�#�� _(��>��n�,��:U����b���O<������6��dZ�d v�n8�A��R֑��)z���cx�A�@�u�@�V��u�\��X������rg1P�֠N�n�0�7�*���&h�mZ�v�Dt����7�J#0d�4*�����H��e��-U2�"�A��+2G x���2�g	�w�H�����cQj�wɏ�8uJЍ���a��3��:"�t <��6���@D����+us�6�}�N��d����&=�����WU����Fz��m�?�1D��'r�ag^���&Rth��C�q\�̆5�H�&�w��,�a[�T2�}��D�5�� yd���Z����s����!���R�Gt��i�,��5�㴮>�א�=WU��x�ӽ�О�������K������H�҂�V/ff�
e�	�Z�8>C���B�<c�;�5҂���A5oE������jtnCh�Hn�;����7"�@4D�|�du����V�SJ'E��qߖ"R%�SL�+{��l�z�X��2a'�79����p�tuܨqv&�}ʖF?�t��KQ5�����M���Nd�9��Z1�d��FiJl��t���aKD�?�r�q�L {�Q-U�k@,
��^�1~�ƁRt8" o�$!��7�ǪXs}��K*q�$�!��su��9�n��i�a���2�	���-��B*>��P��K�7qdYS���@5Ll<�<�� ���8c/kI�U'᪺٫Hm�Ѩ8GEY+~�]�xL�ݹ6ɉ	��ƍj�N����e3�|l��r,sGF��/��d�v�"$����Ĺ��+
w*����S�O;��
aIZ��������|}���}�˅bD�6�����\h'i�����(^U����\*-���w��&��<l������-m��5�����%���C��b�t�:�{��é�ԑ��h�*�����؊D2���X�6>�&CR�E��^�XoӄIІf�%��$>����q�q�
�&>f
A�l����_�D�v$� %s	& �tK=�6/tc=�p��XȠ\9�������Ip�. V#�1sr�y��l�;~�^��l�&��r�+���*�Lk"���q��Z�Z�I�ekW�5cΓ����\�m̒�>B{>h��9|��n�h�߳ÄQ�@�X�<�!(�����}V|E�vS�������4�sX��b��M�m.[�Լ���v^�R��&C��kAZ��$V�\P';�X�, ���%Tٜ��*�����V&�_wz���#��,7���zp7e�zc��(>���+�q,Va%��1�ʚh/Uմ�l+��B���o~j��ם/B� �4��nݷ�G&K�)��UA��sJ���5�V�}��	dq/�i��("5~ޗ=a���k��b�,-۵S`3H��tF����4�rG�.݈�K��	�^	�<����\�c����>#|M0W��0�K��OTc��q�%�50}�ڿ��Ҁݍ�u���pw'�
�N���ji$���ӡeHm�ko�j7\�q�
����j�;|�u�Ϛ�/׍ks��<�%w�Pb!ʬ�����j,F��;��;�s���f	P�E�-��6���J-bmk;[`h��'4(>By!�ņ%��� ��#����S;�����-*v	�] 0u�+���Ų�S��c݀���.�BE��D�V�Da%��N��A@���[Msq�I�H�}Y����}��Y	h�#����]�$���C�a�Q�[1��c��z<0��� ��P�q��a�4����Dߎ܅Ax�"=ux�W%��"X�V�w�$w�=���܈��)}3
�q*���C�?<���L!r]ӊ��cC�KP�lg�{ħ�J�B��<���gA�eȎ��x�n\�pYf��������'�B%���l2�*q��Aw�rĳ'N����u����	h7�&s-� +P(������81�@��
��=;J�슴��
D�T]]H�2#R�랣N�8�*�7���t5F[� �K�m	��v{��Ј�w({��웜�R��I!b�8m+_����NE����oJ]�;5�`�ߞ�~�"'������s�+�cD
9S�X�����}�u=j�
�f@ �'m<����˃ ��u�q��I2s�e͛<S�z�G���H��f���	�n�v�D,�-{�j�J�bs>]6h�ooÊ��X��Pg��*���F�`O7]�_��$����[�kq���'h@T[�`�t��T�����6���N�$�rko�"�����7E󽹼vQ�z��e��u�.��iq��y��0����҉(�|�Z�(3�G���z
GtV���Y�z����K^,:'ڶ5�mge��p�n=��6��MY�-q�w��rW�ht�������r�nZ�8N��<�c����=�����7]�N�`��`�� A����l�/3Vݔ�����q�h�ޫ7h�9��8�d8Ib�hG�3��	?4#lL�/	�V�����r�F3���N�ia�I��6��5q�J�Z`~�GW�7�u��=GWXe�N`���2_.~� �<�N7�v�&�m���a�3������PQ�<����ؘ6	�B�߲V�̣�bG3�eC��	=R��T�[����ԟ)L�:�)/O���F0�3�)	�sz��r%M��z�=R^h���.�D�(�m.�ṉ�|����G�,c��彞iw+�?K6l.�>�3$s����&~OF>�	Ħ���_��G�I�?k�Ø��L��6���e �e�����q9� �(EW�t��2-�L��\=���iw3[mrgג���"E�ر����]ہԚ�`�de���n�\6�$����b�H�o<���S��
��F���h���ܺ;�+�XQc飇��F�R��_�w�/h�[%X�M����6Fm�H�x����88��vx�EP|4)����!,!.����������3z�XԞ�bJ#Huz���#�$�l^	�xFa._A7v��6�p2Y�B��w�h�v�"t��l�#Tw)��#<L�����N��r��'F=��f�P�����g b��W�W�5�Z�v��G�=}�f��QA��ԙ�Tf?�����+J ����z�����.���O�`bBu�th9?�������p�;�9!�r�?����� �~�_�����ˆ��[����8�޷�V`�a~|Ϲq��.���<����&U/36��诘�
�������.���:{rY�qlr�s������/�z���蒻�`#�o��{Z�
�/kL,@���Ϭ<�Y�LyM|��3�f�5�x���z�Tg_��Gd���]KZ��+�b5j�{���vSu�GbH"�v�aG��x�a������4������]1���N. n���$.ҩ~�^k:h�i+���,�:�E*k2!����k�[͒���q���MD��_�q:HU���6��:b�s�?\���Z�m��V�|M+�����ȉ���Yg��u�^_{�IPU��vK�H,��l�A;��V�����ڈ�����������R�"\D�H�y� �?�c�Gv�Hn�X<`��G0�����$��8�?��������-�˅?K�^Qq���W�v�	;qZ��q=�2�/Ֆ���UP�m���D��;pN��i��o�D:�(~�)W�#V/���]�r~�X'W/�Q�7��0�[�j4�d��Y������m�[.��|O�ݏ�}�n�=�C����/�(�i��}����2�ʻ\�X��y�I��S��b^��X5~���͂ej��B����%\B�����XX��KB�]�C�w:�0�ڼ7��qk��~��S�[-{�٧�W��b�yfh1�5�%f���6L��o��x�)s���'F�d��ONc�<�^_z���7�$%���SJ]�"����8�:0�}L}%��ؒ;�z�(�XZJf��Ж�A�U���h0���&��zC���4�i�[��捶ɀZ|[s�;W.�R܇��:Z�Z�"�n�q�!��r��[j��⋡���;���4e�5��҂@|�k�S��\�!,/Ψ�k��4ݯ�
rՔ� �՚���7����		��8'g@e� ���v�wV�=ȭ�=����Ɖ��|�\�̪&+W�J�`�f7�2��P	���1��v�$�t����!Im ��_��r��,�֣����a������RWyy	)<����N@���l������vX�N(�":E��ǰ!q��L�0.9f�3�rn:���7�&�gTF_�+���Ѽ��P�R����NV��N^kL�p�{�W��������̪y�xf25ֲk��.�h}ƲH���2#_�{�ǯ��ze�i0����7�W��&��{���@8�%�a��(7�3����]�Zv�óf�A��@�{��sg�x��v��I���G���!�J�Lۗ�zy�h&>������3Ӫbo��]X*D��Q`��}Z�|�W�v����!`b�-��}�x3�Ҡ�9yX�OL�� f�����v�<}�W�i���͸j���w�W5q�Yb�)�f������*��D[�L
oT:�?1H5�ʐ	-��C������qNƊZ��jC�I�į�N�<#�M��h��?�f�}�#-̗�X�1)H
����OOt��m�p�3?5r��W�!�+�%�7�<.tS�Z�hL�Nxp�M2#n�h���$I<qF��QyǷ�p~�A�{�Ћ^��_�SO�g�h:�$���eޱ�t�s�[?0�-?(4'q�������pL=��y '��ಃ�,�l�O�j(� ]�{B�V%_�p>!��8o����	�c[��YR\�u���`�@5�#�#�ʫ� qF=B��6��K�EW��V�4{
pP�pyJX��q\Y��0�V�r�n��k.������-�g!�?N
��2�(�3ȅw���{,ke�t�Q����K����'�/ΈQ�H����Y/w)"+I!љZ�����9�'�P����F�8@2�y�3���T�JuvO$=J<����ˁ�M��)��:�]�-Ww����TR��"�}��x�����;&@F��㥔��|i%xO�B����%��Fn��˵E�n�wĜ-,�����¿��|�24�D��������ٓ�>DU-��
`72t���Yi��ۣ����M�����Ϫ����ds���᫕_�Π4�j�WQ��Hj�0�(5�z�u�џ���"ғH_�ELYY������;���O�
�!5<z�Ӂ��?1b��?Ċ3Ѵ���N�Fk�6�P�֟���r֢�		^�Ø�~5�*��8�K&��Sb}9 -վlD��};vp���7��л�v����v�!pDVQ�2��u��#��d9طm=F�<2�K�E�R�Z�qr�g-���+cevtR ic��J�*b[!���u4�c,����۝�y���DM���saW9Bݔ�E���:��z��Zd�(�7xd��~"��`L17���4ж}u�/=�`���>�}���,e��l?P�F���+�!;����C��h�(?��+��>°��� Ĝ�fxk+8� �V��.�e�=�P�v��[t'��8[�"G�oJC��t9Ld2��>��N걩> �j���u���]�D<����$V�zx馬�
���EX�P��ᡗ"�w�w��O�����lb������u* ��.�|�6~툳m�"E��M��M���/���L�<c��8?:���#��������咵懄>����:�xe8\�Mm$@^-UDa�c�R��*��zʟ�h+#U.���s�Wˏ��3$��a7�eM}�2+��٢])�3��(�c;-t^0��fc�*�+Ķp)w�R
����u'-D��R��`��6�Ϧ@��i���dȤƍA�]?Gs�����$�f|[$��(Kr�f��c���ZF
�\��"bJ+�y��<-�W*R�#ʲc��Ƀ�r	�q�8f�Ь�N���F��f�s�HԂ9���n�|2��zU����?SgH��^�Ғ�Y��,Q��c�>�(�8����l0d�=r����q�,�EpW�̝ ��2�P<�YYR$Lf-b/�)��7LN����_	
�J�='�*I�AK"�,Ɠ��51���P:�!�h&4�Z�t�.4��t�U�=��eWlO�/�>��%m/T�c�^��1��Mb$O1Y��T�3=	�p��L y$����Uk������t�(/��L6kĘp!J!��_i���7(�F�B�:�y3o�RH��4���g�4HS�$��^[���8� P+J[=/j(�J��(��F�yR�/:v�,���2<���6@6���W�{d- ���0x���t����Xs�c�Ӧ��;M���cw1yL��� m�'��"��{wo@���[M�M���������x(U/��ط�{oya�zQ@J�����ĔVA�D
�`U��F]�����
���i�� Zx��KQ�`p!��!|��	���<N3ݯ��Y%�{��L�v�G�(J��]����=kMea�;��[��J'bk�TfW<>U�1X0�r�$��
��so2#ߴ<�B"S��q�^�khl�(&pN���C�G� s��rղ����ȗ56�pL�&�P6�a���R}�lygE�.�շB����IV�σc�4��߶��b�s��ѭ�K�0�r����6���S��$YUˢ�֓�U�����[U������� �{+j�?/�R39�I0�(�Mw�s��f}{�Rr 2�x1����z$�p��\}�ʝ{���Ǌ_I@@���tj~����^��}Kzݏ2�?�����_0G���@^90�����nvSA�Wd��&_Uw�S2�9n'b��o�䅺9�RD�"�Ywu��ǀ��Aɶ�~Ac�ׁ��f<1�O�@6/��y���i�Z�a���h%r²L�'���ҏ��5S������+���l�����]C�Ó�����w��K�)|��ű��[�n����^�o�N�ƺ9����:n�8T�2�Hr�s7���z�U?���5��C��u�.�6��[0���� �R��u�ut��q���s�1TQ�Y��j�|\8a]y��:Nc)�&�]�6��x�@�z�DI70%GH������قZH�o�%)�X�j�Z���Ш�ʂ�F���&ZYf��Fp�q5KaX����Jp ���y����P��3���Ւn>�r����)��7��9���&�*L|b�&��)�֣�����Nt3�nc�F��~{{�1e�C�nC���@d}�B��ӌG�Ʌe��w����lT�»�f��S��.M(B����A8T���P�7N�-�~&�Z�gvb$c����MPY8S�6!�;V�p��H��ՏT@]j�qN�]� /��B��+~�U��r�l�I%��*/�K�ϙY����QG��^��IX#̞u���������f�������q�>�+�1,���݋���-�8戧�܃6�J0�x�z6�S.��p}Y/����vo���o؅u� ;�e���c���P�l\N�
��tM��zp�b+�����>+e ���E�p��
�}׶֚M��Ա�[4χ�S������9S����͏� O�/	���S�d�
�2�����G(aX���,��5g���/��B��z�R��cu^�q�զf/�-shA��^[��I�R�^ ��XٳMMm�j��L�%��/�G
"bh�h�	R�Qs��3�^�?����'Ge��R%�b\�"��<�ب����9<���ܿ(t���#��q@.E�ڛ�5�����(�I��gY�@Ӥ2,�Ԓ�Z1L��پOa�Q+R���Nw;�Y6ܨ�U��gI)�� 	��I5��_|X��Wz_�6y{�L֤[�5���du�K>ڔ���2��P�FX��/����_���{��$ڵе���p9��
���Os�1$x6�� ��^��6�����m�	l����٤�W����o�K%��T =�2�\w�@&"8�Q�32��Ds��v�,�c�pĀ6#�>K��2,�K�U�s����%`��\��"xt^;�+6|�w .~t �\&Y�����o��O�B�O*W��|���o����!�6
���������)�rM^��	EX�~�	c�j�Ep.�rwX�o�&���\i��d��#M���٪VV���c���5]���zh�&��£KS�{��FRN;<�I0P�)!�!�B����,>Z�6�~��K�͟>j�P��<5�ukR{U�)b�g����N����%zX�B���q��,�@�&��S��H7�����6��q�z��w8��`��\2��wA'��=A�z X�����'�??�]{E��4�����tL{(?c`�k��JC��u�p^�"��AZ��~��FS���	�-ϒ�E����`)(���)!�Ϡtc��D���o��Kvb�DXlxVHYEB    6184     f80��!�l[����e"d	HZy�e�+7:�+�r�>��3�J_:�i���B۸�`6J[�Jf�
�+Fl~�d�ռ�)aܗ�Ur%K;��$	Y,�x����	�̅�Ϻ?�b�k2�rV�|��]�����D���0IX�"ԍ�B�����c~�^�a�;��X�
��n�hwF�UfvQ(u�s"^bNs��D����a�]ҾW��hn{$��Ǟ�:+ �v���\�
��Vr��`��C=�UO�����D|�CUS=Ha��?X��5��Km�]���k���V}����͟���j�V��|�����M	tZ�h�Xf'���(���G��MY:@b�F%��B�[Csk��a�>�nd�� ��e�hV���ȼ)�!b~aL+t,���P��vόV�-
3�zx_C��I�cjaA�+��?����7���4��CD��9#Qx�^��(x���h��v1:�I�z^~�T���ث�<�^���.Wr;N�S,٧���3���['��C��'Gf/r���H ƽď����A�;uHm���b˖1��zgr1Ɏ��Y��J��Q�T�d �}=��3�>0��UD뽤��Uj�*�	��uz���S���wd�f���d�a��\@7���Y�C��f
��-���F�]����6)��'�z#}לho�3?z^��\�mЪ��Sp�I��99��ÿ<�[�)��v��C�4or-�r6��hs��+q���s�ʯ��A4V���ҥhL�x�l5{�,�B懨p$�
`�ei�z��_�;�W�tg]�!�dٜ����ML��R3��k���a3�O��J:��Dm�>���^jM[��?iβb��.��/�J۝2f��P�H �}G�X3�8:��D�Xс-{?�s��w,,�Ii���nV<�lY�vQ?��N!�x_qNO�j�G_�"����;�H�m�`d�1�HA�?��xD��w]��LH�Y'�Wb,�-����P\I'`E����[�	��� �)��	W��vz�HÉ��ω�;A%[���<Ku���j��O��Y���L���|:�U�0L"�( ��"<����1 ?�X�oo�-���/0���Y��狫�n:Gx�׮�9�q����ф�dH��d[�7�}ѱ��T(r 1M�l���/#��tA�iz
כ���lŒ(+o�X�)F\v��D���:z�������6�O��W�M��Q>ĝ��V���:�U���զ�SY�^�&�2/#����ܱ��r+�� �c�r!�0������V����En����E��J媐1�W<�G׼)��Bf���s9$~�'띦.���W����A�d��ƫ�;�$)B��ƥ����b�`ͦ�Ԥ��2�����_���
�p5!*���BF��΀~��^�U)I�%�
s��Q!dPP�\��٥����f�L�c�/��d�/)���Y�<d���HrV��x��>K������M����ro�cj6l	��nk�D j'E�v��b' ,2i����H�
.�|�j�JX>+2�e;�yO�!ui���^��֡e�(4y,ӭ�(�5$ն�L�Av��m˴��Ã���I�fn8XaR��#}��[��:��4�́��j��ӕA�
/)��:�\2��ё����sqN4�
�]���	Ó���<6�_/��F?������ˇ�S�3�`r���H!D6b���(pfX�6�l�ϝ�z0��4���1Ԑ�XD��գ�cAd�4l���5��Ӂ�h����G��Y���F~�}*�x��B�|+l�t��/�v��,6*�L�v0>����s�I���f�ʖE*dSh>��Ι)IM����~
����OcT��ϩW�, ]L�{,E;뙡�l!|h��jK��e������%�j�U��/��D'Ç�t*B.%�w��/,�7�6�����e>��g���>l.��{0@-���(j�W����Jd�D ��Z�.j�v�஖P�,)l"aS�!Eӽ���r���B���̑m{�b���=Y�J�O��3n�.�ܼ����8���hg�":ˠQ{I��z��o~�����$��Ӱ�T�ы [�T]��䓒�K�(��0�iDE��W�_��M;��7��^6ט��}������/|�U7� � 9��!�&���^�:��%g�y���$�;huB���jC��Ġ��Qt�L!9�;�f��qT�^0�_>a�|��nOI0�OLe��0y�J��s)��}it�%����"�yh� ���|H�͆���*1����oL��´�.%U�:B�y	�Vc�CfcE'�f��ؚ�D��B�7s�n,Pa�������.�"�*c��
����Z`C���9�زċCd��ª���Z���7���t���� ��z�f!��a�y�{E�v.¶���0BE�a+kw�Ӱ�Pߟ��J��c�]�:�܇�\��k�yv�k*����h���4�f1�����E{$x ��%��}N�}$L}0ߛ��ᮘ���Ls��%���!wG1bJ�`+F�")_#H��[*O����6��Q�����(H�!z4ڥ	�>m�J�z
���M#��J��5��v8߾5d��t�#E��~�J>���u������,"�BgA��U⪛I�.-�6�7D��Md����Ԛ%\��v�y�cFfZ�[UՖo��#"u��qxHZ��wm
'8�K�aI��x�⻆� ���"�kG�	K�v�����%���$yMʽz��\@D+<.��� ���+ϩ��+E�j��������9�����M6�ij���U�~�ˆ>ı�d� ��";f.u]�������Cϩ�J�`_���E�1���ȇ T���b4J_�ktP I���+o�(w��FΒq�Mb�}4���(ˢȘ�$�[��BK���(9AAc�Y���^��W^n�>1�65ќ�O�A�a�,eC��MKx��c���'|Tm�U���4p
z_d;��r+�+K�d_9D�}54�`�����V[�����>BqȴAkwӧ�9�G��	�7�Zkj7t��`���"��ՙ|u���H5�1x�~����aI9�Y�L���D%����9Ck��@"���Uҫ>���H�s15X�������J�i��?8������i9�P<k��X��"I��Y�\n�U4]�w{��ؖ��i"�Du���]}�F@-�̩��^"N��t�l�Z�SUK0J�l�O�-��k^����x>���6X��#Q����k=a���	>��eD\�m�����j��g�k��ķ�bwed������7�h�YA�`[�<��(� Nr��j�{�O�����k�O�q,އUX;TT���T��l"Ll~<�a��$M}�����!�˳� ]�|�Ք�'�������!L���l2���p*�����
qW�������N�l�V�~YsSQ����s$Pл���t�U6;�w��Qb��z��p���מb{����-в���f��j��t�����ߥ_$�Wyd�%y���,%����wh���k8LJ)9�3ChG�{��.y_�����S�GFO�P��҈jS/_%�sΉ(o|�JuӢ���U�^V	}�Y��|��u�ڦ�����}����/_2�sm��� �+�h�$�w��9�$ɪ�;���~��� B���<q�;#Al� A�5�̳�¶e&P���K�?��a Y��o�%O�PƋʙ��팴>@��Pa����������X���q�ϮCU1`�6�kl�`r�:i�!(1|v����V�4�]��7��yR��e||E"�p}��sz��	GY�j����U�*, |ÌJҠ8���:���3�E+'~1>��N����lB�w"�|~E3�Ø�XK$���En�����bK�C�������s���