XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��2�C�e{�k�;�*=O�*v�	�W�A�b�����.e��sB����Ѐa���Y7�����s�2ŷg�݋�6om���F���Z.�?�2{�!��+G�I��O�TV�B����1�o*�=aߤ�,�M��7"����Y�cO���DN�z:'j/��_Ү�=@��1�;���a��DG`�%�S�t���v&4���F���M�B!L=��u�y����^�S��H)
�#���y~V���q�̑l�M�A���H��ӧ�����H��uNa�?Ò�i�Y36��<5�!<©~t|�4p��ݔ�4�f�m�l��ᚵ��9(E��D3Oms����<W���)'�J�-@]�I�ʱ��@���39�Ҕ~t�K�2�T-"$��u5dhw��@���Y���#M��8��q�2�W���@F}��˸�T���ɏ���ť�M�+o��v
@�n�JviL7���ƚw]`�K}�ѡ�ZU��L�6��͗X�)p�h*ͨ;�YT��MJs��0� �!�[�(f蹷�t@�²�*M$ �#�Z
��&�m��>`B�@q���a�S<�8��ЛY!H%�*�J��Q��KGD��/@�[ ���0Y��k���~����p5��w(s����6(R�&��K��F��	}�9��}��Ծ�$Q���ʨz��R��1�w1�u9��������n���X�XG ���i���ڡ2�1NVF3W@�u{?6���R�(�o���W����Q'#n������V6XlxVHYEB    5df6    1510����iC�;���uS�������8�U>���,�H�Q�I*��7��d�C�'�}(�5�8�.��z����96KN�G)�}u�c��η����<�/I?�ܸz�#x, �uI=|��+���o���B�I$`�@a���羹z���/�W��Y���rr���m&�d��a���sw�"�7�%��{;����}�]�e8���K8].xCՖ
e�:�X�jQ�JYc����vg��,AE���J�섐��K��qȒ�s��h�u����lch��>Jc�#����X�u��"�77)h5�va|nm�}ە�^J(�OeF��~�Ƣ�LJ�zJ�=���x�-�8 �� �|�C��#��\Mx���D|�m�OǄ�orŎR� ���Ĕ����2���'X�t!������*�
��� ;�R_�#]oJ���n��o��rV�aF��/j����yTĩ\�
���Xġ����D�e#U�m�����m�X�io1�v��r�+0V
��r�_��h��������˭�&jtG���~��3��WR�rR�H��Gc=�ڀg��#^���={{= �Bu����~1��t	��g5�@s��%�w�x:r�<D;�@��'Q�C% @`#6G���qV��_"nl���V ]r-��~a�����(�=��?7�o����L������:|3������qTXS��+T�����Ψİ���0�_�B�m�w~�e�@�{U�C`��Q��9�M�28����T/q�����b80ĝZϔ,!)�9�bfAm&����nWU�޷��{��3p@�b�����5�\B��Բ�����i��
W�:�8?uˆ��!H�5!�w��:�>sِ�`G��~�HW*�'�d7O��nrՁ����xYN17�abX�r���7_Y�X��5^�����6� ѭ% �k��4刑�c� S��)l�c����be�+d�bdV��m�Ė-�I��7i�I����{��Cӗ'� ���q���V��?:�!xVEy�v~`^�uIR��M%vIף����߇���T��y-�j�
���!̂2��Q߼���^>�ҵ����yL�[�?�v�����4��T��L�}��WC�a�U�F�y��Y����!k5�^m��H=�dl�y?���Q�Ne�I��<����ߧ��1��n^ї�
��K'I�'���m+c�\��?�W���ؙ� x�/�w��^��z<ұˇf�}K�<UA�k�W��A���Л�812G6Y�
��n�#�O�au��s�%�J��j#�U�%�9�&M��(����q��3�?pOOhV�E����qL%��IC�Z��9'-�������7�{eȐC�v�+A�'|�Qϯ
���g�� ��~�tT���1�I)�����gxA�-�eQ�ǡ�LEL�Ux�ő��u���ne�i�w���աP�ϴ�9�l�˷L3��Ֆ�p4�X)��}��0���{��6��AC �	�V��0#�H��κί֏gi�G��L���ѤE��S�P|����5��`��s��ʁ�.�����{��</K�$�'&"c���'��������y�����"̘[/~8����+�N�k�.�����ZJ� ���� ؆�!)�!J
�[�O� ɳ��N�M���X�^��w�Ҁ���@h�j��s�68��π�&9��o��J��AzW0���h�M�DZ ��Z'l� k(�FIt*O> afݘ�*���
z;,�۳���z@4��ɤ����#�ك�f�%�0��Pl���ۍ�G��2�[S�I��s��m���!|}EJa�<��X3o�/Ѫ�]y��,�U���b���R�X�Phzz�5�n�N�aE2K�K6���Y��$i[���	�w�2�����pk#)�g�\��9�O@V������g#r�\������6�-�ƍ=0w} �ZJ:��^���q�#�o�1���˖L���g�k$�E�r�tM�7NG-|��N��<�7��^��
j~�#=8��1�k%ݣ�,��Xٱ	;�;I�����e���;���3��=��D�$���gj��P}���(s����-Kj��D#��VFqX	��i7�U���[Q��w^�R�=���up���~�qd5�� �	�|5�GoZI@��'qYl� ��;�vOr�kO���o$�ޑ`�W��1�M�#f���lj��aD=Fi�ئk�hB�L���4�?�Pd+âq{����Wr�#�/�����l�
Z�+SC��y��R�m���h�_�P�.���ߚ�%/��J�����6�T�qB�7��(�E��P���R�iv�>�O��l�Yo���(�ɜ��½k�����[)
)C��E�;�_�>�Rl^�T3�sTsH���8�(k�gH�+�������ػNgX׭T���-��8.j�B�GX��z������Y��^�ݝ���3��6�t�<��A�u��c�BY�L�ܶ���z8�=��.����ǈ���!�5�>J�R���)Q`&$��<Ff�k�
��|�`�@��ɐZ��a�dn�w��#@�Uъ��k0��JT�ӉWe�Nr_�\�R!�M��$�r7rc7��]���mK6�ڗ[�%��I��g�UVy��8���� /��bZ�Z��˜6�Cn��ew2A��RG����Y�̇.�$Y�/�i�j�O���7��c��&��k	��J�z?ؚrB�{�p���CPsnȌ�W����t��t<5��J��>]	9J�f}{wϊ�S/��V�pf�W�t�XR3�t��rbR-�b����_�eq����
�#��������]��4s�������!H9�,j���k�nCƆ�������e^���!d���|��(�GWZ,��)L|y[G��p���?�����w0 ��{�b,�~�=�n��T ��$5�מ�ؗ>�|������� ]�t�L�Κ�֏�:&�<,YB��e�Iw��'�ª� ��z�c�8h����'��hzJ��n��7�����%�)y���_ �k ��3h�}L�N�G�.��g��3���V4E��x�,u��E��G�mz	�Q�"��*?��M�`U�k�#�H��_�q������"��~|V�������4�	�$��Hg��W�զر`9o�f���1q�`UB���%��X�F���:��+A /�¶���f�����J�)]n$l�$���ZG�MBժ��]lWR|�)\{ۍo\Q�K	�T6;������<�:k�D���*?���I-��QsUQ[(�R�o�2�U�nG�	�Db�u���m�M���(>YҰ���u�uQy�2�t���%ʇ:��qﴡ�P����HC�.C�R�.z�+���ق�v�R��@��H&E��1򰌱�3l����s�1�%~�)_�����]�Y�ӲJ�Il���#�[݅E��%�l㺅�eعn�qyyϱ~򜒶)�#[W��@�1#JV���C4��h�mFeJ\ɂ�yLJ��n��*��N�)ΥE6�;�8�x �ю���?}�t�aI"]��N�6<�T~�t���2���D�٥m��;to����������� �xٳ��Y���:~��92I�/���v��&-d�ŏ��]Dl�>��篙�����Zx�N��!�4�>Y�Ydu��/KH���'��� �z�$gf�k��%,.�R.��
���ϧ0��)V�G�?��F�K���_�D�ڦ���yL���ZN���]홃Z�_�l����7�<�=m-��}gg-�m��,����4
�b��y����8���hv�W-U�ho�(�rB~�ubJ�0��\���g��PY���{���2V��T�ɜ;��MQ�S��n~�A���D�&%�xj��4��:M��k
��;�\�r�(�����A8�����OƓx��(���:��
�H��f�^mW�-��fh�j��m?��2��N�f i���@��YQ|>��G�Ւ(J�{$k����s�:[> �T�L�,�q�i��E�h{���h[�zU��xw ג��
�_���f��Jh�,�#O.o/��t�c*Kt�ܵT(��,�ݤ���.v�c6/[f^GA-h5v �4��z����Y1��ƚ�m���o��U�Y��Fχ�a���!�y����dU��ƺ�4W�Q`=�ٵ�Wʢ�Eо�����/���(�mtX���5�g���|bzW�7L`а�Ք��s眭er����k�%%`�[�峀^�>mk��P��f�X�%����qm�/��f4���b�7�� �T���P�j*�5�� �=x�;��(�I��ð.�O���qip	 J�֧C���F��-)rJ9��(�|_/U"^�xߦ��63���A>��k5o,v,�i�U�?�ßB����k6�M��NF���ܪũ^���B�F�N����O'���0Ka���A��	Շ˿<4��=cY����-�ծ@+!li�+4x�h(�o�|��࣍�[�z��Q�?W�yݦ�z�ݞ�(�t:�j�⋷�FsǪ�˚�9��ݽb���a�s��2:W��b��c���3��L�F�½8	Naߪ�eMr4�6�߰�`O�s{�N��_��!���pD�Mk6�]��cD9�Udd���y���
26�]]J�ޏ�%1��$4&�%����w�5�nF�,?���/;2��7fs�)OD�T��tRVlX�0c��<��o*WS�j3[״"��ލgpe򹭰Z����Lfl<��|M�jБ��
���7C�TM�Bir�M1 X.�#w��PF�e��]������	�	"(�#�	S�$W�3 ��>�`�5�y���c��F�by��֢o�kX#�y�`�&���ʴ��0�ACXwZ���F %�֕dj���O�!z���Į�S+�	@|���Zs^������$��'%�qt׷A�\ĭ"7�Y�]�I���mp�m� �j�|�ʈ7�7!{�d[Y��{o��ֿ����b����9�����i��n�5ǣ���9�C�E��)��U%�G�ݴ4�z���f�5_=|J%<��������4&gc��7\c��_��$���aS�wgo�,�mў�)�PUv�?��]�T�.`M�v|�7��#������N*}ۢ�}�ڶ����5�,�:q9�Q�d�|��֘;�Vʒm���-q_�E�D �~k~Z��V���x��*�l�{��Ǩ{J��6g=�E�3a�2,����p����%�v��F���3a����