XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���9J���!���WV��X4��f�"�}|٩�8}�LU>�kc�s%o�g~�w|}
�!�vW�O��p��M:��T��Ʌ���ZZ�X?�?~(�,����j�I�U��H��!��E@��y+�G�]O׉Plf1!����#�O��~�G-j����3�<`x�����_��;ԑ� �m��̫� �T��:�_��gJ����+�0H:3�4_,�����a�Hd�F_�@>b�&�J�&��S�(q'_�X��Mz����)�#��{�ܹA��n:�> �D�R�[�ӒtJsrC��oTq+������j;+i�
a⁤��F;��~���7�a�~���rې����(��N�(�R�3� .�&� "+��q��$�. Հ)���m��`��'i���,��R0t��'Jj�"��U��z`ҡ��NP��:}?S�Ǿ|]�����2��"S��"����^��o[ȍ�j�)�7�/����g6�ۉ�u�S��$�`�G���>y���8���o���x�lCϔ��w�J�Xg�����߷\�r#+�M�^y$ѓ �Ϫ�Z�ܚSәzPo|�# }��o�I*9V~{D�dύ9
e�K.A�[)������N�yz-��2��I[���
Y����Q><��[��U�Z��X���Kd��ʹ�f�	���F:��.���ť@_RY)�~`�����o���|���{vk\N�6��a�#���ߤ�/)�Ԙp�yQ�O��Vj����ccqXlxVHYEB    761e    1770%���G!h�bupo<��	��&��9E����]���v@�*�N�
�L]H�ٚ�3�� ��}���7%~��Ѕ���X蟋GV�D#;�>��Ƙ[��H	�(k���G$�����|��:�^,7��fދ��m�T?�QT�nq$&�v�=9!����>f���q��s3Wʾ��:�L�Zc�Ĥ��BG_���I����p�npo��EI�K*҂�����&��MaH�:�B{<[�q_K�����C�S����T�-G�����dP�?�gE��r��+s�6Ǿ8k9���=��)����D3�2`��>ܖ3O�{r-�fҢ�dV)�KD�-���"ީ�.�@^���Ȓ�d����wnP�Vg`�-8t�&_��[e���xtJ���Ey��WQ�p��o����Y�²�QYU0\�	U��)h����n�Te��k�$�`'t�uU��z�Q�gm�a�䄩����x�����-�J1X׶c�)�ʑ�p]��" e�>�||������)(Z�5��œ�T8������.]�cJ�2�1�-/
�l�&����I�
[�|��S�׶���q�ޥ^%*4��O<!8�J��������K�xۮ�[�!��&"�!�A���i׻(,g`���'���{A֗Q��"������%=�~ݞ��� �(�ļ�^�IT�vEy.Dg=E`��*V�_�ԁ���QOr@p���G=h8�%�?�X4�����$-��~�Y~n#�Ծ��(zۢ� �*�9!�9�n��Ƙ�"������s������
�,Sm\L�w��IҊ(=��T1 XN�Qr ��qo��eӦ�M���^:�l�y<���P��X�`e���W�!s�Tڷ��EHš��1U��M��[���{?����|�3E��\���_"��@�52�:#����$��{�ɨG9�q�"��"�N`e�̟��1>�~a��
�
�c��9E����f$���܏�T��U:���ͺ+&D�\� ����<�7x$��`Klꊁ�k�'��s*=J!�)��4U��:��״o&�9��yh����zMSK<��mI��֨kZ?�9x���e0�.��^���տG�2O��ɔ������$9$�Z�����:i��2�/�A�햼Fe��8G��O���n<�UɅܟL7�7��*A�(}��ջ��F"٫���/{�dq�Y�q��1E8�F��!�+֨�^m��h|L!*�JH�B����$F��5���*~��M�#^�Z��F+��6r��o�`	!Ge��T��晗��F��=
KA��]x{G�.�ڤ������4��HOkEM&�?iP�'x���D����0�7��ٳI��`^ t��i�5�n��P����QC4D J�O�HXON%�ba�_����/�z�mt6�o8�e�����L>G"\���u'	I��㈾��-��M.�{fa��"��^��T<�9�- nk��B��嵅3���b�]�������>��^�H93%S⓭������kۏ���l(���S�д�ڂ�ٿ@��P��o�Ͼ�Ūq6{��I�3���Q9���܄ُ��4���:Eg�hHF���̿r��Tn�ǥh��~��n�j4`k�}ө{���?&�������M�g��4��0m�2P��f;sE�"CBw�E�	�~Xf<�r�U.��_dl%���`��s\���_�~NX�������}��O(�i3N��~'�x3�^kA�&���	�5�4B�@�
���L[I�58>��BF�bj�w����T�ꍔ��-�d@\__AJj/�IAN.�,uZ���c_�6�BM�Ο�Q{�wT�D�vF²���'�#{�����O���'l�ji�FĠw ��4Q<$i۟ b���{� �*�ܒ\E-AX;���X�c��6�n�2�aѨJ��n�k��䊵��f'԰��<0m6
jI�7��
�R,�)���p�@o��.$��1���S��k`?����f�=��n��L�+k��)�}7�r������noS��P�)�v�W(
F=�����Ws�k���P�3'��7Z>^vt������4�tS��	����5+�l���I��(�+�Em�VuHƑ�")�l��� �&����d��5bcYc��U:����^�y�
k�v�Y����l�lc��~�̰�}�}�+tg��T:@3l����j?��G�nM
�
���ʣ�Yt��XF��c���	�-�9l��B�㧊�;d�n�s+hH�v׮���q*l�n�|&���پug������K��	8l��i�_$ͻ�aȌ�v�)
a�LX�e��]�CjL��3]��\�q��7?NR�JNR�[��#d�di��qV!"K@0�h�#�e��\Y6�������G$��g���[0�$ jw�b��Y&W�����`xO�&��Aܫ�Q�$���JpO �uct�QlӔXuRL�R c���~Jm�Y�J�sn��Rc���J�����pY<���V�4`%�a�_��̥�V1��Xx�N2g-`]���|��)�i~��`Ϛ0�V0�o�<G�,o_�_���v^�ǹ�;��\��������ܿ���nf����/�U��g��_ϝ'���]@L���\?:xo/�%3�9J�¸�S1�G�|7}����`P�<X89��5�c���G�y��N��v<����-�b�@*�_Rl�3��gǽ�[L|�z��a2,����K9���G�@��������Cc�|PY1a������Y9Br4u�����w�?3j��*�]�wޢ�QP���jD9�ka'� x׭W�c]U�$���
k����P9���,R4����@U&���J  )6?ڏuM �J�&�U�^��9=���?��yY���B@�{Ns1qM�t�1GdE��&�5P���9�FY��ik�=$�@;~>k� /C}R�c��$�VpNj�P��� �n�U॒��5�YfF�8s�p�:ܫ$O�~'�b^]M>�����V3���@�b�z�o�`7!�҄�=�_&�}�V�1ò�>
�<�9�8�Y�ᲀ��Њ<L�w}a u�@�KQ84���7��؈9K�����ո�;��!�i����T��r���!��'��LD���툳�6�H�t��C@P�&m��Z/;����aCi
4��/q뾈�%�d��T�\5飼�˸�U�����P5	�<�BكP,�߮F{�n�^8]�!!KGc~���X�.k�U�4]����}��K�Ik'6Z�l�,���x�7��1��]����m��������vXpMT3�J�4 �7�	�d��3^��w<O��8�y�������ᣌ2��(�����D���{���:�;�{���yRs_C���/aW�b��[%�kϪ�f��>���k�q�"]cx��m�	5i�4nn� �1�e_�{g�|��o<�g+��@7��4�"]��&��'�ǅߨM5Cr�{�� ���}ok�w�����ױ��&&�����`T^������U�ʹ�%�|m�`1��!1Ø(_砎��6-�@`$Kx��f��oX��'
�=����z����7�IC�	��Cx�k����������,L���O�"�ĈG��4�#���! ���^u�k�A����>�O��� y׬ۃ�AG�3��lj�;ī�zΉ~��B��f� �[�Y3�E��X~[�	�MbcJ��ϝ�T��Y?�j�,��\�\��2�P�b�����/>�9�8=�-������p�!j��H��NЦSTA�˝�Q�Oq��`^+��,�:E�d�Z.�k�?�eM�o@��^α��M����zb�q奼?(�N~�\�o@�K��?4�g����,	G������A��>�����q)���ml�`��xD�e��lt���)�~����� ���f)�	eM��LX��O@�L �r�T�jұ���P���Z\R�8d~���-+R��m�S�jy�mm��k����N
f)�ԹQȭ������0
|G*<{���L��E��� R��π��\Iơ���ͣy�Zu;�"�h%��|B�l��~�V%-g$�8J�}*�̈́���OPk�$L�y�)T���̰S Ԍu��Ź�qBBi��Pb
�2oX����a�:�|�\���ɣCGȓs��s������nIã׷�`S����mp��$b6��|E���ȺJ?}U���R#�g�	y?+V�*b����Ze]>rE�C��I��d���rYzK�5P�B>20�o�f7xB���c��ƈ���ϙ���E֦���bm��'�a�h�#֫f����X�>�*ԡ@[&ܸN޵ԿiN3�3䦩Lo�,��yQ+	G�dթ��.XD{�粜�k��P~���px��؋�VP3Y:a�}ǫ�mK�QaZ�ߤ\��Ro��q����R��;������!�_�}#�|�?�0���] �9upp�g�-�-���q�bT:�E�sQ G�D#�B=�ll-��'�A�N'�u����_6Y_�g�`��	�D�M���U���C���|A���n��}�c�����e���7>2"���&�L�c��!.x_.��V �U��y<��8�7�MR4ѡE#�j�d6rL^��tT����;$�>�О|�}�B�^C��E�Z��+$��i��-�����@�E���P��E���U���|��y,Ll���L��*D�b�1�b~�_��5��\��u�.�B�n�!&!v���Ř4�X��Ѐ:1k�DT�A���0�,f�_f��$�Z�j�`z�ץ�xO�x�:�r2Ј��S�[��y�P���,�I_�'!ۻ�7��mOt��{��QO5���MIA=�	O���L?���'ǌ6eYF���4��GV1s��T�I�A�ޝ�Kx�"��@�7s~��P1r���p|=�И4�y�'j8Q���S�v*K� �
�Z�*�ML��2ʔ����-$��P-�oַQ�zq��p53F�+����������$0�nu��ʑv�f.��(�l��l�"��	���V|�O�<Kj��&&8����:7�xE2�+�����û��f��$<N�C�"4 ����1?��@��؉4u����^M����X���΁��:�v<~~y����g:��w�d��۲�| NO���\f���p����,���c�n�3�34�M�{���;K�4�7Gc�E�Q@�햳'{���{-���������VL����F\�2���}��i�OE �u�:�5�o�a7�&�ٌX�1�k�4y[*:�ni��g��#��@���%��Lۃs�S2~>M�J; �I���RK�A���0!QٗYC��f�J4;��i!1���v�NTO�5��^�9������gM����h�7]�^��Ojy8�e-����1�������jR���'&���DK����IL� �������\���ő�C����1���	(v{oI+�c�e��4��~���6'�=�
�K�I��g<š�e����cF6ڔ�BBE��8�2[d�����yF�DmAdE�}�''�m���ҽ�+�֏ ���1K��ȍ���k�u~�Oo�l9K2��ծޔF%J���<Q�+�C���HAmh%��U7'�a�u��W:IM��� T�&�����B.�Nt�"?B�5-�5�uС��BIAKR�1�↟1h�479�O+����X��[:��$;*��$��~ �P��Ȱ�yo�;爘��-@o�������8��X�{�a���7č�wv��xv�Z0��k9��0�q����

�����7�e�3n��n�,��K{)��j�-Y�M�ӵn_��TE5�E��H��^Qo�}p�^�$���7�S�p���eY�� ɳ�����e T������̍\�d�ϼI�1
�@