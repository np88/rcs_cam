XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��c��AHM���xx�|	6'���?_*?���KC%}�_��^�&����n�/�; �s�hs�'ĺ��s��sz��T�#J0z+�Ήu�ގ'8u3�^�����AH�峘�A�'�m�[��ι��׽$v�X��]0y"m����V���4j�g!M;����f�j��<�0�e���4�ԏAD{�s8.�2̇л�j�,���� -�II��UJ,�����0�@-`�3�����_�(�gM�;�o����9`٬&��i� ��p��r�š��)�W�$���\<��ʹ��s6e{�j/�x�d��)��qʹ��w�IzK[!��g1�k�H�oe�󦑭�֠�go�j�w$>i�9��[&H�6�q
4�\�^�����GU d�Qܶ������#"�����m�S�"���A
�!����z �E� �Yx��w<a��y_g�0��[�]���Bx>�)��_����j�2u�c4���UW3��6�`�'�T��:�D�0'j�JJg^�o������䧱[눏�^��m�щ'�a���'[�8);�V�m�u� �ȲvEZ(=k|��2�|�r|�?���0� ��oL��$ϧ�=,�nشB�I_����Gk�]�Ӹ
��2�:���iqo_��i\r��{K&�n�c��*�R��!�Y9r�v�E^p���=M[���ZJ�os{����C��h�ȕkzFo~����l$��M�LB�S	;���M;O�h�R/��-xԪziw��XlxVHYEB    7744    1780K#Y��i�A5\��"
�A@2�+/�#�>��&�7��pS��(���� Yp��e{R��ĕ�7N��J���[{���h���O����?k*ו���6����u(�� 퓨Uc�x纼�o����-��~�7a������X�����.���L�xv+�G��d��}�F�I��f�y�@�A��RD:�"�6>�(����� WV�Bj>�
��t���Sv��~0�Q�?掠f�CbFg@,�	��I�軒S�����-��|���W��{�fUA������2��p��a���i28-�T�(�%^�l���nY�'�VΥ�<�h����U�+�@e2�7e�z�l�7��E��姱�=k-��� �gMu�/ix|��c\�9��{nW3²�&{�s��v��δ�ʠN1b3�RK��������N��*۩�a��	��dA�Ԑ��q�^�����Lw6��X�++�s\Ro��<����������ʆvA��lW�!(ټ����[���s���>�Uy�Ɨ��.�Ѹ��_> v �dQ�n]w3���S���1-�U�d��Ků[��o|r6��"諊%Pe�����[�xi%p�i�[Qq����c� �r�i]�s�0�F���m�t�2���Ma'd��̪��!.�#n�b���l���0(sr�$�G�H�n��)�C	��I?�\1�v��>Fc��Ӷ�㳔5S�#����Ȍ��!s ͺ/�Z5�2sD?\h"b#=�7KY��;n��(إˢk�����R��]R�Ǝd���jfM�	{��`�\!Ͼxa+(���|]����SYuk�/ۄ�?�XD١��?��Y��X��c	�R#ݜ�������������0fػ�JʼD���Q�;s���-eR*p�Q(_�~�����,�G��v~ p����0�%���8���ſ �2��+�\|�ҕ��.;!�	c��`ؖ��B�`+�a��ה�^�p���'DA�/#��-�a�V��1Gdmd�	��	B�%�`��jKH-X����C��Q��/�s"3w����[/S{�P�����x1it��r,�k��v�|�I2FW#>cukԺ"�Ñ�U�^�(��ݜ�I�}7_�k���D<RX��+^D�x����JCAnY���&�%iSG����>��$%�w1=�H�Y�ѐ����uz���)����r$�B��_����H^����3~D䤸a�Wi0���w��兎-�.U����ڿJp5�̓����敠�9�(?'�����,[�ߥ��/�':l���ԥ	���c�Ui���J�0���(���\�DS@����~5���pǑ'����5F���
(����ٶs�,GL�p�OK��p��1�[Tk����e���~ ̓�U?���o�ϯ���;�`	��`("��?�:�r��r�����ӟU�V����^+'=o�kP/�N�	ΕO�W�^�j�#��B"n�bt�����"��/w��2ǀ<��	������ܐ�z�u<�x9|�Og���$!9f�qMyI�s.!MT�?�E��DKM'7����\����i�i�5���lg�I��3����N�o�ٞ�y�ekKV��� ���fF��Դ��� ��i�\a(�^ce��ޯ�_�鞄�1:��|��kY�f@**�_<�[jt�@�.K%2�"^�q��&�OI�K�� B{S:Lޮ���=����|�2_��aZ��24���;w�[�f"a����O�.H��Q�}�a��G��zR58~C������}��6���'p� v�BDr�h���j_V���-m�W�5$d��ΌE������㙛�j9&F��ΘC�*��P�E�ʨO�6�Ā~���&��_]N�})��ʺ�lL�L$e��H����҈ ��$g�E�ao\s�å��ie��t�x�=���=�z����8��hf�r)�U��)�,��U~�ؙ�u���f*��[ٝ�P�}��H4��yS/-�P��aD���h�?0����GmB��X�*�H\�ɔrr1��0X�b���:�2�{��M�ɚӪ�i��p��$�HҴ�fڽ�^�?�^-:�-=c�G�랠~�l�xw8����~1���	0-�&j
E��8�v�7]MC]�M<(/~3ǵ2vl魢S�9��i�3e��=�&*	^��0��J�F4(;�g/%,�DF���.k�E�s���ł�Q!
���67Y��bj�0|n�_8	���HH a����җ��=�B�m$⾅�U�5����J*lӔ�q��uM� 'Ȋ�Râ�����9�ݿ��f|���4Czm�-��?�M�o+�!�L�c��V3�������'rT���KOֱE���?��3��Kp�j�O{/ճA#�,E-���
�Ao�={�]��R��տC��Y�z��$U`���K�ë�R�Uw�$�h)�4�%��j[��񓿤v��Z9�v,��u���#Wq����P}־���\ ���_�5 ϙ�P[d�?�cX�)f�J�U�1���)Zy 벵��.�W�Yf��>6A����KēV/!�}Ʉ���5#._$����c�O�ct����6�2$�=�י�t^���0HL��qʙ'����^��\%�b>�K@�������H�
0 _��1V)���¤h.�`��TO�'}�R"���?��p��I�P�`ps��h��|��5\Z��[ ��dǚ�y�9⬋�l�K_���X�7�v���~����wt�XJ���
#)[T������y��a
��Ip �9m-2�z��ꔫ��l�����Z #���&g�W���Rpj�J�<z3�GZ����7���5ґx��j� _�sB�^g'[M!��8�M~=�寧����\�?�s4Tkovz��j��$�*x{y�n�G��/v�&"�4�I�lXpc�䴿���n��H^����f�f
�+�@���@nt-���v�>�|��Ӕ�r��ѥ�9Ìx�{l�Aw����o&3�U,�kd1��ϜϩZ����� Kz�}PY��LKG��8��@1�J[5�qT/܃	��Z>�D+K�Bl���U�S���&K٦eB�)�=��������Uh���0��@A&b�hD��y-}v�u���-�&X��a(M���8y�lv��NB����0%4�۽�$�z�«�#�6��6CiW�_*��g��(��Y1N��3�Ea������8�{˷�����P�����]﯉�y���K�F�V������h{��2��e(��h��1 A ���>	$ӛ�j���9k�ʠgX�,��3K��I~jcp�g��#��ŕ���
,g��b��������g�pe���0Ӹ��`���: �C��/�S+$m�,/��kĆ�,�)���&U�>����<U{X�1��1���Q�����Sk�Bϥ�] �����p�L�M[�1Ҭ��b�Tyi0Pl}�e�i_��:b�P'�A�"1�5�2y�Bg�l�j���r�(�s���Rs��雦�4x'L�W-B�O7�yذFS��6��Mt,�|�Y�v������P1�l�%0:9���k�<{��
�qn����x���Qd�P�5(�q��!��-�-�v(�g,1��e�yE�" VNUK����R�p�p&�t(F�[,�����h��N��,�	ĳ��D�/���D.��(gk��f�kK�ƾ�g��w �����c��(W�[��y�Eo L�m�p ���P�͆)����4�a̳�o<�O�6��@�_�"#XM�AM�lP)��8�C���S�U���3�/	>�f>I8�{�q��99MQ�sG��ߌ{�"����QG ������Lg��b��Մ.��P%KDh�� �7����Qa�`�gD���ς�U��g�l��(����=�0�
Hg{˾�#b�s�50�>ݫ,�|w
���^w�R��Q�#��+���f�ȰJ~㏧�I�z����E#ͷ*�;۳��M����~0�����4c�pZ���+��2�PR� o�G������ż��NKA�8�G��j�n�:t@�c;�,SZ�5�������}˚�2Gfvg�����ʶ:�7U�p<A�yL�{ 0+���BD��>L�m�	q{�54�`@J���/�-88�=��NpI>������� �}`��X՚���<��c���0���[Öͷ�,�L3�s�[������5��w����0�h��JPEKU�}ԑ�z����2��؏$xc��P������/�a�`볞��q �y�� ��jn�E��p)a�N���zL��z;�ƍ�����?��ױd�"r,sˏ)֞g����W�c�񆥤���E�a/!����#g�T��@ik�;�2|��=z΁��&�w���Ѡy`ո:�c�G�ùd�K�i�+�����G3pۆ��r����+$&��x��)Z�A?jv��A)���X��ɍ,u�Gy��L,r[ũ�Jj�QK�����>en��Zg1l7A��u��*`��T���]�U�P�n�/�d�ޝ�(#Dߧ�ɪV�����|>�Ņ�6X�F�(��S��&���^�3y�$�I�����W�s+ےV�����
ܩw~A�h5�ȸ�щ���"?i]H�	oC��~0P���ug�\��o���?yP��7��.��l��$�����S�_w��I�5��r�;y\��j����6�T�H����Γ"S)�7c&t���P���Ӫ�*�J9����-���a�V�ڂ�̓�zb]�i3�+zRSn�&i������ҡ�a ��#<ZҀ�ߖ�9Y	%��@�Ȯ�#ϋF1��U5kI~d�������O�ꕉU�0�4S�>�S��
V��_gj�4�>�O���aזU��F�u��?�'��Ur��6��k/�7����Z�]����2��J��)	ASܓ�ܨ�Ud���m��2�@GD㜷�р-ly�ɥ�ҝ�kx9R8�8�䙫ݮ��K��H�p|W��+W�5Ҷ�}�%p�s�1���Y�S[�ܞ1E,`��	.���6Ҹ�"�j����)b��v;�a6c��
�ЩX{���6�m��Ϗ"�t����LJ]�ҭ`�F�3���Џ�`�3��,��Ux���]�,H��M���o
v���yZ�:�at-{Վ�ܞ�|T�:45{=�n+;.�Qks_;VFPb�T�<�<߾�Q��4Gx�3�x?,��~�N��'�(��?�N�O� |u�1m���>��v>
�#<�i����,pJ�G�9����*Հ�_�׽���f�f��v���=���˩����{�(�ߟ��jvj�ݸ�ӌ�L��{��L:����%7־��{������2����A7�j������Ш;�`��w�K�x�r�l	��]��4����|�ʜ��2,j>�0��M;@(��$��e�(�d��[�挍x
T3��`�#��e���W�W%��nUHI�k(�����ji����>��G<T�]���	v��3��;�����yev�K�G)���� @!�y�1�|���rMv���Մ���~������)Z�{sV��l[�8e�֥e�1��ɦ���M�vm�9A?��y�!��H݂�\����F$t�<7���:=a��С���Ǥ��~���_3&9⳯eQt����!�~ ]f蘷;�KY��s�����xZ9;������&9k N�?�?�A�Ũ�:���4���[k9��c�'�+;g����\(����.m�/�d#a�Md��{��85�18l�n>e�$ȣ�=��+x&���S���>�q����m���hkI�w}�
*,���3y��5��׽��T�����Q�yn�b	� ZL�M�)AǱx���-�P�5�}y�=$���v��F��1�$QY�