XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���z|
���7�[Fzk�{�L�,`�+*�:�Ǘ�
�9��T���������)�����=���]ZL�LA��I	��C\\
�l����=ß�V��%�x��(�����.sg�����)l:�RH�f�qF�Ǽ�`8k|.f��&V,|$j�!)^�y9 �w<$�:Qc��y-����^k����B�աf�Ľ9j)�V�0�(���+�؊mt��u{	ЯK��P��J�&_/�`��,�!\�q���]�ص,w��P>W.N�4��5k���9�p����_K%<B��D�2�I�vR�ǹ}��F��e|����9��g��I�'��\^�Di����$L/�[��la��cU5�zZ��J�.xhE�P[�9M�&��V���Gʀ��g���Z1J~����IB&�Dr�k�ٍ�x^��w(���y�M= 8N���9�0'LhS���.U]���`Ƕ\n��Aԡc��+(J�H���`��	��{���,�$�q���{F�w�7*�Zl���E��U2�g��ga�[��	)\�>�z�I��>���/�[L=�.��t�m�3W:G��l44�
�J���P^��7���JJ�6À�I(�k٫�'4�������m��|��b�Cw[��kX�C72�t$:a7�-�����g$���dU����|�nG���)EH%��=�{5���Їn%��=��F����ݱ�SP�.�	�CUNˁU6#�5+����`�����""��r�A��^� �/�$��=�XlxVHYEB    3504     ca0��{��(g�
0��D�׃�nvD,(.��mR{�j���HAW�פ�\O��ʾ�+� X����'�[�;�S�F?�xY�v�c{�.z�J�&��iɩl���Wƌ�F��6�� ����$S�d���Ϸ�<���9�������zC�R����`{�����0|+z/c�6��;W��A�&���,?��/��s(I���Z�!`j|:M�c�e��(�͌�r0�(�f�l��l�n-���r�g����[}RV� �����4�/9��3]���|�yk��S#����Js
�XV[p��P[d׎f�>=��+wĈ�N��큩�! ����oQM�]�+VF��5�-ށ��%��I}�g� "֚,��M���.?���g!R��o t������"��`Y0�ϵ���q�\fB&��?&7��}W�]i�O�4�Xϰ�{)ȓr��h%�]+�p\�>���-"6k�$y!����>%E��P�`;Ւ\�G�W���'FߝX�I�_��-��jĠ .�m�Z,,5���a�/8��	#��Ra��:^�{6xԳԨ��jĭ�C����.�O�&@s��r��� ����4�
*kF0Q�=���o�b$���8
���w�JM㎱z=�R�ů��jك����Ф_�]`����v�9d��(�����N�J��Wa|=
'|	:,3�a/�J��YR@�PY��lɍ$X�k4r��)��g��1�M�,&���v*�p�p���:���ӄdUTtQ,���}�x�-&���icd�T{ Y_lcYZ��^իa+\�U3��%<���� z�6~m�,*L�Ҏ[c�@��͟�癦09F��\�\2��'�hċ[Ԯ��[yd�a4n�J'ƚ��������7�̛7m�/p5�����!��"�,�P�,���X�Q�[(E6q	*�U�'��M��%`k��6nP�� �2��>�/KZ��h����^�8�q������yS�Dl��hK�g�l�_ڪ�Z�a����FJ���K{��8��?�T�&�G�.�`�*6�q'x�i1_�dE�sbp�Q����(i��;�o�~Pc�[�tpw�u�n�Bo�p�ą<��O�d>R���}>�S:���)c�����	�>M�7�%�����e����Z9;�3��:�r��֥@�Ҋ��ȃ��!8A6��	�D8�"�6�cn&"��UNY~&���e,��섡�,Oi�"���B�/��d�|�n�)�.0�����3���x�vp֖�[���j��a�9U�E��(V��O^���~A�Ό���M���{T~�O��̣�gruBG���;>Vif��l��2}��``������n���rK�7أ��t�3y�T}N���*�S�����,��v\Jcxf5�*�ö������aZ� ���QX/{��:ks���Ds��7U��%,�Y;?:pR\��x7�ڮ�O�J�:W���EJ�B6�ym��sӇ���כ���J��W(|�N&�'��@�-�TG 14��5�<AaP.���9���CX�0��<�Dts�a���"����L%�e���8à������������UO�P���$@�5�Oa9���Ȃ�vnF�?Z��Hڮ��+m���Ƚ�K\��&@qwa�dx9�j�T�?�,͎e�#GT��X�ZˈGF�"�/|����ak?NM��L:}�:fB_6�@HfI�m�ɥ����E�~��n�+�
P�N!F�����A���d��5�$�Cs>��e��M<���2)���58�'��N��Ғ�^�x��� �u�xo1#�������Sяv�z_�^:KWU��Apn������b)v�3�=˂��:Ϯ�]�����z�<9�'���s�����6�]6M�s4#���������B��^���5���������*�j[ȥN����\�G���byhL�n/��A0c����R����F���;���o�nS�v�D]��D:_� ���Ew��] �Iۃn���;��)T��:�Է�O�E﷐�;|���O	��y!�9���(��%��J�e��$ny��xhH�m��sŎ�^�!+E�]��^;�����Q��z2I�̘�+��0C,%�v/Y�}��Y�M
�f{�/wJ���<��*9k?��2zn)70�B�I脩���앧F�]��>0u�,��xL+�{��]d�[PU\�,��`ܘ=
��R���+}4���Cа¾i��06_� ��".�v��ry�����}����N E�l��b�O��Iģ�M�䑢A���5�iqF_�W����TH0ؔ��ϧ8����N$�uX�J��Op.(������oOY�D��>�F��k��I���HB�K�ʮ?H��=.�,'5z����D��p�#4�(��8�H-,�c�=	F��(1�pK�z*��b��dh� |���Ș�u���}���F���\�-��Ø�h�����$�5� u6���RC�b����/�+i_,D��Q��G�1����@g�}�X�`G�i��I����%��1�4��=���ΈҶ?�_��o�5�
|����P/}"/��9U��>�4��ckMc�٭��1/�8oY��f��*�:�0J
-c��C�G�e��QIL7����S|���'2>)HYt�`kʻ-���姴(h)������%��q����#:�sZ�]�Vd�L������]����%�jJ��Mp��y��G3&Ooh�EZJ��o�k��P�B��}�4��1}�%r!�N횓���)�M��L�sey�����	��]FZd���N�����(���/�-o�M,Coȵ�d�vB�t��ـ�]�-����L���������RS�_SH��@�l���2s>�~{��E�k}�Cg>ʹd�j�P��2+a�M/����Ȉ#��z0�M��>�����e�)2A��l-_�!.���.�A������ad|�b��������������!�Qz��f�`�zlE��⥌�^�u+U�4�����+I��LQj��'�ux�9g:���t��t��O9h��F��Zxʾ�~�lC�f<4+�L��s��4��"�zh�z׹B^׾E!I	9-YT[��|�.����@˧s�4�f�(H46kA��m�0B�!k2i�"��