XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���N�v�Z'�5��
��KI/���29-F&7�Z�2CC���w#�hh;��R6`b�oFf����	�n�-�E|�U_�GA�ǹ:K��3k�#�D����̲��o�	/0��[�s�j|���U��)rA	6%K����&X�0 v���}��a���ur���B�l�IR=�\/r�����u|u�˻J�#8jQ+�Z���y���`u�!{�~�V���ہj��J��IP\`6(y�r��x:�p�Jꕠ�Tr?^AL��<Y��1�x��
��V�wn\�O�0PT�K:���m.i�h�oBy��i
�3^ܲ-5:��P�Bp�e���iFpSP���Nh֜>[���VV��T2��p�nn݀�Z�A')�ѐ��p39� �v�q�צ�(�������G�����mIf�����˨_��8�K�4sї�*�d��Njz�ӷ:�ZW���Ԟ��b���ͯJ��M�u�ѳqv��Ϛ#�׫�ˡi�h|�9+U�]���C�\	$�	|�<����>4�	/�����\	�����|�A�>O�)�0���t�0;�\L!�W����e��b�%�gU��h�Hs��A{�Es��2Sw�
��âiɀ%ݥ.{�r���<����"ՠ�9kw��Q8�$��'j���0��Գ�;n�RyɁ�x���0��Ӹ�I�*�$x{8ޮ����Z�$�&�R��(� �����<)ٵKvp�����X�RG����e��TXlxVHYEB    b380    1930�u`g!�R�3q5$V�vVo�T��eL���W%��H���z2c�UɈ1�L�sx�ʋy'0Ƙ��3�;���~����V(�˕���1�T&���h�P`�5���{�����.���Q�2D.Vm��B}g9��&��~�*;�K�����J]�Au~VA�#��Y�V�Spź����ă�X-~h I�r��l�B���Iu��;BE�KmW�‱�;;�ܷ����D	���N�ڱ�
5T�!��Ӫ�;
y��Z�|�x�x���44}v��?��9������/�mJ���dx�6*r��9�ꞁ��$�5^�I���a�n�#!��h����bs�5���><M�?3-B���1+�M!�HXf}�j;��[�����ud7/�R��ԽiwU���L��J�d7�� B5X������j��76�(S1�T�4���.��=�f�}Z��n�B��tI�d7�ėT�駕���l��r�*��3ik{o�ȯ��-���l��_u֜+���!7?�"K#<9���y��Gs�qS�|7#�sx�:9��8W��~���Jg�tzM�8O�=��i��?����V2tw5���MU�)VvD�K!�}�ߑ�7GУA����`�aym����tm����[��l
2!|�E�����p*�O�e��ʛ(7<� �A>@���*1�1�����K_t�kr�9��c��c��C��?O��BW�0�)k���o�R5�6�<7�Ô���w�ge�܏UU��<i!����|��w�Qc@���YL����Z��>L������3?QU彇�6zb2Y�]OV���>�C�d?ʵ�"�V��*�(jRw�q&���҃H���\0l���+�2E+v�A��K�b�>ȷt�cf�6�̩y��((x5xu��w��_C�,��]����	P8�K�s���$�SܷXg�2L����L�3~�fo��BB'�	���0 n&�
�.'�H����}~{�:���l�+���g�A`�0׍D���$= ���y��c~����]����A���k�qaI���ٷ�G�1��@���LtƦ��Q���˥�~h=��q�s�7t4�wm�����7�ͻi��%o�)xf��N;�/��fy>߉��{G�s,�������߁��l��M@wޚ���
��!�]���D��i=�Qu{�f��;��b�Y<3hd0��Yg�Q䂂����!MIF�kf���V��&�������|�S���;�OB�/x�V)B �Ә��Ͼ����pv��dq���7�
G��L'�I��Ҧ�~8Z��d�<�K���0��ry}υ �������3�R����{��o��@��QXu�E(|O?.i��#d�X�F>�p��yf!��٠�գ;Ws� �׆a�83�P�+D�����y�z)�o!�"X}.7�����^�k������R_�2��s�2~v����n7��c�m�#2�ײ�B��.�����%�$�(�R��h-׹�8�ˋ�4���?F���Ď������l�_�|�9��E�
�ǽ�E�ڪ|mSj�E�%�8��
i�hR�.�_Y[��B�Fi:��r����Y�	�~��۔�7�����?p��޾��|�Xz�\]�8�ȿ{�74˥F;ґb4����v�z��΅!�S5O��hƮ�i.�A�>E�kcP�/�+��l�I.������0kJ�tċ�g!�JmCV��S�-jS�Q���[��� [���dX5��9��޶ѿ"��j�I�b�d�JD^�;���T]�0-�B���pH<T�1لs�)��V$����ߺ��@���oCB|*��e�'.m#|�6�#Aq���ԉ^�ᝥ�%䆪���	y#�Q�Kx�4��V�޹�	��r
�[S�H��7b8��g�XEn�g�l)�w�$6T:/N/maFD�mk��L��%e�pA�m��[���Y���I�c|�FҀs��b���pHXU(a~CB_#�F���~J���U��P^�\�AdÊ@tP]H8W��y�P��Y*�j��,O�4=�?��+z�xk��Se)�5^��R號e��h-�wL s��n��s
�y�E.Tw� !B�$]
Z�V�y:�����Z��p��3������l�r��y���V����pk#���Z�ם�m3}�zs��L9�-�]QM���-�sYܣ����mS'�MF��U���ӡ�J���6 ӕ���V�E�x$=�/LDi�0��Y
*�O�f��-��GY�Me��3�{��	�Y:&`�cl�?c|��M�B}z�ǵh���;�0�*|��82��5!15E�*�H�����ˎ#�>�l�.�NN�<ZO<����s��Sm@nm��>��ZH/�c�3�B׌�'�6S_L0_C0d��:�NnHpI�?��Urh�G����#8�4�� �zY�G_\K$����7�F���[~i��H�������Ƿdzm�G���0�5��)u@g�;��e�P��Js��i$�7�����w��2~��BFf�ŝ��B��Ǳ2�R/�O�0ဏk��%�f�ۢʌ퓧۴�m*�1e�n���:fJƱ�2�Ks1_�
4y5ғ��9!�����]TkF�T+��Ք�c�__`�wҖ�b�~}�� hn š1�m@��)��Eag,�!%³~͛�R����O�.����54j
vu�nD��K�j�kR�~�qɯh#Y�`C��r�^Х�1&˪��5�ܚ)�u.��K�{'^y���9kz�L$�3T��A}����6O)�,w��}$�s����ٓ����*�j ���yj�Rq�{���d�X��m~ȏ��@`��σ]�S����[��'~_�� [�%�U�&Ȕ븹l"���>P����.#C7�OL�C�t'��,��_��Ƶ�0�:���!�˿c:O<��*�\Ѥ� �9�9K�ey,]���R��/�L��X���T��zB otV�i"b�j���`�<��Lあ&oB�\qxm��b4)]���׃�S޷c�������f�.7��%����-n����o�E#�}�.遌za���Ɓ� ux.�R��5.z!��n�F�����,����S����b$$��r �k���Mfs\զT����Ej��k�MbR4�\��ǋ Z@�p�b���k/m��/]QtsRs�-�`���S+g�nt�;"�$)�RH+��mB� =�����!�o���A-�-����\'�<�M=���gزS!ggL�+�b�lx��E�D�92�|fK������e��_������=:li�z~C���O�
R�l':̲���'������[�v�{R[&!6vCȜ�N��#C׃��{q���.�-��?
���i)�y�>Ç���f��_{���&0�y&rFOC�.#ګ^V�b����6���:��T�j�v����!K���{aiև/4l�8��[�D�JO4:�	j+ 6�؄8}qc���0��Yuy��I�
��E^�����+k�O��,N�y;��U΢Q�����lC�SIIJ�Y$�^��8�����8�������@��[�P0�V����=�<�h���
�u�%ߗU���N\{��8�m��#ƶ��}7�`g�1�������i]I@rҜǤѕ��,!�������X�_�k�`6fS����a�Ի�r��&�����(%$��A3�3��w*V�!9�k�w�Y���4�^��a�sN���<�D��4?~U
`/���3%T�*uR�4Q:0b��9��E��, dюhrR�"��[Yg�%��ĳ���k�M�<Z39�ь�˵ԥ �&��$���g�g*��Ƴ���Ԥ{}|�_�`���A�ݔ�|��6gM1%����D��z����'�F�P)
Ԉ��}�*8��1zA.ea��,>= �aS�V���j.���K���Ś� n1س��m��?��
����!P�U�B"��sc�`ǥ��{oA�&&�~�����:x�m�D|?�VrI��˕c�f|ց��5'!t�
���ڬ�҆�W��O�E<2@Ĕ���?� *��
��'�W��D�g�(ZU��+~�>���p3��]�C�jzѓ���k�2�q��D�*���7S`��:՜m(����"h�$c�M�)�v?E;���|��c�j;�^�<�xQ&:S���Oj�"���q���p��ꚥ�aC��R%����+ks�����1wOp�����������C����/�����Ǿ%�{�%����ȻbC��F�´E���U�,������^Xr���y9P��֪�p�$BQ�OP"n�����C��W�a�}21��7s]2���
��	i��o�`)F�N��S'��F�f$���7��J(�SU�F��m�3�U1��N%����>��^6��wʬ�I�Z�]�x;��A��Nc\bט�O �8D"�s��TPL�ڑ��b��eA�4o����(Y�N�7pB�ӑ�J�J�jU��f<W��LMc�������}��Van�~��Zt��������x��Ĳ۪�t�.P���y�l��W>���`�d��f��7�h��T�6Pw��[�\�rX�ʋE�;`�6Ё>�ʜ�}��%�(n{�<w�@6\�fi�\��F*k1gU2���J�W]�h�~��\�̖���uq���ӝ"�^�V>3������a���	�ʹ�Y�rG��Rv\[ƯI����)���CC1�j����^c+P��|6�)ýV}!�!��&F. �y��GWa�.����O������LS��U��f��ƍ�ߑ�z1B��m��p�%�[�ز��gl���S���,�iw�a�D<��I*h����M6�dD)�C�� 88�\��}?���
��;�C�'I��c�<�>���
+?�������$�gSŰ����i�5ah547_XqЛ������aA�� y���^ӯ\a�܂�*��B��h���I!2�o��&�Rm������$���E΍�Bp/���	;k��-	�w2�kҤo�^�Z���\ m��u��9 �92V.��um�Y�F���] S�h$��[Tk8�T͍d:�V)�cʃe�;�/WA�L�G'{`�j�ϝx��D�=��X�QPD�Aj��h�+H�e��E&7�j�隯��%0s�������苴l`�O������^ayH��$Y0���5s�.e@D��ʀu�'@M��;jJ���]B�E�m�9�`owĘ���r�8U@���p�zw+�`�/�� ������)�-	ˈx�K�Q����x[
�:"f�Z/M�-}BL���e!���v��1�@E���'������Z��RGc����J�(��U�5�ڜ��
�: ��E���P +*�f��%���#B@�vN^�pQ��F{�c�-�4��L�A��'w�VO��81�����?�ڄ;7a}nc����t8<��O�Cܠ��uP���%ZP[ t�p<�@����/�*��1C�~�!��g��}�Yt���L��?�Ʉ�6п�0:�@�@5��A`���I�b�Z����nN����?�|m�� �j�m�����B}BK��Dx"����:T�*Xo-k>�(��pۭ^"=,�$���q��|��ic�.A	� Q��J��/�k���J�����7|s�hX(G�R�xeQH��m�;��@e|°ig��i)��j����^�v���Ҭm>�S8�O���� Ld�
Z�BM� �{�����l!��Vm#���{<kt�N��㒹&+��ƒa�8�!l��o�p�j�]N׶)x�q@�rT�(�w ���W��DHD[��� '��Ќ��^�CsK�t<;�Rr*����#�xk�V�p� :BH`3���j����GNJũ]�j�EO<x�/]	v3a��A!��a@|?G$��Q���]\�����#*f�i�y��H@>7I!_�� Z�+��r��C����n���>A4sc����=*%��[4����ѿ�݁��@�~'_ُ�3��wg�AWԆ���ȜhX�{�S��lu�X���97��q�[�d��+6���(
%{�&����\�����J.�j�%Ik���N(��N	�:<���揻��x����g����r�3h2�>@jp�Q�-�+x#�݂�AFL��m���U��9�F���-���U�q����+^�I�Y{�g�u��Q#}�2�bwA_!>�5�-�G��ؖ_D�96�-����ڏ* �Y*�L0��-t�'u� ���2�I����l�<��_p��-uK�>9� ��D9���B-R�IGʀ���x34��&�=ټ�'���[�����f�3T���|��>�=E����@λ:�