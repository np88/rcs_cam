XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��[_o�CR��W��θ��]/����|���ki���\��f�d#�Kx�[x���q�G/�Q�[�Ul�48y��$�`�����"�����j
��Q�Z�\� #�����v�rѼ�gyG��M�\8���8��l#��E�k28�l�_�~a��fI*]n9Bٓ7���_��)<U����$@�&�K���QH��sAg�L��Ϥ��9�����v9�H&��}�{?+��u�����I�3=鎾��չ	�;?b2EI�s�ߘ�t�
-��X����
tGnf=��*2jӕ6�z�ns��PoA�Fv�,�Lg֐�B��������Q7��17�ElDW�U �_-���(,�i��+�	��*~=��x�k�9����(��h��ր�K�ԡ�C�t�K �L&�q&�	���JH���µ��xknۤ�/� �z�7��ԭ�U�'?�G��q��4x4=�ס )2x�
�Y��d&ګ@�k���|`pU^�.�#]�#��5)��X��� Ln����b�T��������	�k(=��m���Uz���h(��*�I�)1`�^�/�i<���6�]�"9|{����o��&��du�V9�Y�X�H��S#��@��x��Ol'ы���m�.;���~X��0��^�|��^ڢ@0=�n��[_�`e����tS�v�oZqhV~Xp|~qI>���<Hb�,v�G�C�F�!z;��.��yZ����H�@5u�~ϛ~>��ʝ�Q�/�/�S�^R�mmE�W� \�̎�0N,�XlxVHYEB    55a7     e50M���#]'��7��d�c&t8���ٰP�R���3�v������/�p��u��XZ��}�#�,1.��`G]f�5�./�T�K��H�Q���[<j�� �F�����NT�F������N�B �S=j���"�8+D��"cʝ&8�T�R���T�ԑ�<�w�i+��cӐܨ�M���L}^7B�La��	4-��������� ���K��qţ�$�۲7�x�_RU��u��h3CM$Iś���"��gp}��������s/S��0=61R9�uXtz�qv�q.̸�Y���,���zfu���;0��H���o]#7���n}�rubG��!m���ʷL)q�H�c��.���DЌ�rn����6�
f����#��O�6҃`mfǗdՈ��8�}�6�[�̿��<q��Q�0�8-�V��v1���m���Q~�zK�L���d;?^뤁,�ԴDC}/ߏ�u�� ��a� �U�D@�^'ZuU�� �#��-��h��!5Q�d$~}�r��T�����ɺ|���r�0���6����	�u]�_��؋���r���#�[�n��Қ\���L��M��5T����h�J����t��'ke��f��0d���+o��θ�O�,�`��Ӫ��m��H0/�9��!�+�[�^1�N�r�}&>;�+���2�h��8#V���� {#�ҝ
A����LWH�4��Bh1�JC��M��@\�L�O���G�GZ�H���[�&�]�d�o�a�ʚzIK7��`���;K��������::���w���cwV ��W/�>�U'*����	�[d�'�P� ��,�,���C�ю�N[����a1|;��o��X�����̟����byoI\ʈkc�]Z���ǭ�g$����.��>j��&�i��z�Y\��?:���N'�[^�z�g�ؖݹ1�c�� ��*�!�\�*
�������`����+#�z�;�tӊ�"ʣ�}�"K�3T��de�Σ3���gz�����"�<�U>�ѡ~ϰvvދ![�u�}��3w}�����0�V'�`G��[�a_,ΐ���������������� ��R����;���L���U�6�Od�6O(�H,R���������}6�$��iҌN�����E9g�@!�:�!0˓>ӛ��=&3(��6����[�dϨ�9l�5�w�ä��m��L�j�>�_q�[{M;~��apJ�n�X���]�خV0O%����y���,n����e)�ŞNt����ØZ?�t�u�>�r)XѼ�u��,&S~��W����Rz��^/����W��I����d�V�`�ca2�)�k0�7�#{�w*�ᵽ f��3���:Jm1=[�4���� �ջMP`l{��ۡGa��4�K�
(I J���#pgi�Ig\�C�i�o��l�g�<��`����Dam�9MjQ6h�I�3��B�=�AJ�����)
��ٹ]��߀��*llӘc�ʟ�8-���E��d	����{������00yn����-�<�.�'h��!�)��~JŠ��|�.F�6�s�M�Vh����}ݧ���L��?��W�F�¢��-��N�EtN	|og�2i�Q4\�ڇ �ߎA-Y���EXerӞY>�6���.+���oY�c�	��Ay���_�� T_F Ӎ�桬�[s!ɏ�T�?�}ki�B���
(��h���K������f�ަ击,�EB�Mvs��)b^���I�&·/��������A�v�MAK��-�Y˶�(ߵN>�x�/BSиƃ~k��r܄j�yC�"X�I�`5�}���s�U$�F%y�V=�Uz����������<�i�(��'�$Y��D�u�(��[
�a��"�GHa �<�}΍�yAbb_�=ED,Ȝ �%��v﫸7#2�&`E,C&� J��;.��nS�R?R�u�P^�Y|;ڸ\R	���MOڎn4�!�0<D�ݴC(t��`0��N��J�//
�䋓	 �h��w�*�3���^�J`^�	�ٷ8S	w��p�-ہFz$I�(5[��T�}�Ӵv5�������	1����p�~��@7��������5�K_�,�:Ӥ���Z|L�΁���YB@�����s����~(^�Yb�8�%Y�i�-�M$S"]#v������?�X��Hm��8�{��d�1���6��d
��%�+lA��_c��;���Q^�0�oi��RF��F�A����f�4)q-��_ ���A�n���K��`�z���\<{���� y����L����*-���ȸ�+Q6 �,�ɒ���6u�"�E�0��H�fm#�B�uu�<]��_���o��Z �᚛rt��E'j������P�a �_�����=FM��!CIȔC��?��4-o�15��»EbB�O�s��/_?�Pm�zDb`zo6�xB�q��K��*	�9���DPa3�Z�*�/�������	�j|���]�dj)�;J�xfl
No >����s�[�����`f�{}��?�`�@b�!��J���خQ���Q��c��uc�h��GX�s�' s���#���G �>�CR
� ��s���6�u�M��a*�cُK��r͙��*���S�B�iG5�=�J�Ɣ4c Uf)<�m�̠��3���c<��M)/�������K_��:������s7�e�aI坻��z�^x���<5�ش���}�]�����C��e����q��|��f��VZ�W �<��d�C��i��3`T�e��W����l h2��7�g>/�L:M�P��G\j�H�.��B��}��2�(���ˑV�x`�33 /�Y�?r����q�3t;�H��P讨���?#�B�<V��t �ˑךm���\ʏ�?.����ط��ޛy���P�r��2��&�����&��5[-��7�����`Y�� T���H@�6J�Fѹ�ʖy��F%L�Ąq2 �̄� ����D����/����r���'-�!.�S_�U  �L��zj~G���LkĈT+�a���Hl����It�n/��5valw�Y>��tg�������O���E���de:�Ȼ�Nz�y�M�v[;@�k��)�(��z:E�WV��k�T�A�\jz��h �.�_n^��;T������}�9V��O#
�S�ӏ���r�l@��u<��
dZ���wgKn��|�8�E��No٧� ���H�ߋp#9�A:oe�&��TVf��OKmok�����T6��#q���cu�f�Q�֚�zǢT��D�[{xx|$9��܄�+Z��Dj��3�U9����p�?���f	b R�����{���W���zLtz��_��f)�h���mY���	5k/���I���	��$Iy�*%��m�#q?��
*rܟn�K*۶��G*o�a��F�K8H+���/���>У���<Wf�чp�"��;{L4��I�������u�p;2`(V,�|V��"r�k����,L.t&y�Q�^�]���p��I�d�P�zwe�<0bBA��%�6��lc�$P	x��݂<�W��˼���@>�0�n��'JT��#�fh�