XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������#�p%�Fz�����T�cn�}T�~���[��M�XJ���A�2Q̭��*Y5����v�J��\Y`��<�m��(P3�΅B��n�;d�i:S}F7d?,��������&�66Nz�����rڍ���yU��A�~�`+�m��B#g�8ԃ/��2�tO=$�9�ٮ�l�Nħ�'?2~��B��ѽN����+�� b{)U?��KaR���K3�NE��	U2��A��b_!�t	K47�65�D�O�k=:hX���fbK�3뫸���7���J������t�홍��Hr&�]���fE����P�7� �����z��N�L�g4-rp���=���L;�9��l������`P�����������5?_IE�{�y;vLh �X��PA#��0��qJ�bQ�b�)r�G�:���{3+���7��5T}�rU?c��8ng{�f뎻h��S����g$�朡�Y8�e��z�9kb�}�����1��9��V��6pŋ&����Ɇ>�Fu_"�۶M, bjk��7�!fɐ����K�E̜F C�8�+��:Y#&HzޗҘ�����7�X�f� �B^�R�X %�֩,|q�Hl~���Jޝ�ڀ�0�CjڌV_;Op�1s��Z+�S��:�ғ��$�9�dnZ?,��Gu]F�Kى��8�W�y�(�ч���ç7����9�A��(5ze���lk�D���j�ND�h)=��);e��(~fji�!8bO6�"����XlxVHYEB    fa00    2d70��P��֮}�]KPx�$D�}{{#�G���
��?���J���[c��}[Ko���!��a��'g�XP"M�²�����K�?w�N�Q
SXXZ��"�xY$�z��f)��}μ��X��zj��tG�.}oag�]o�k(B��_���۱X���w��Ya��������5�JR,yf�P	͋��i���ew��&�z�z��88B���Z�&��%#���<ټ�� ��N2S��w�r4$�ti:�!Cv `�ns��{�o؋ی��R����_E�!.�Zk�C��FM?y?�|��ov/S�zf����4y]�Tػ�R
v������Z��H�����!jO���ȟ��>%�1��%a�VGD���i=�A��<�'4ҙNO%����vb��~��hi�N1��z;OX)`��lm�m܅���Mbl��,s����Kݼ�&�]��ť�\�
ѹ�+�]�+e��âo��,˻����7��qg�M��ˍ�������{�=��foy��ծ(9K��x��(m�>h�2�'َ��.�IɩBe��`f���To�sG������z��;N���G�%�kb����f��k6��)}��፳3���v����ŲY�m�>͢���Ph:�q9��g�mB���b`��?�y�!���uj��?�-5�}��Bi)ξCi?G` �)I��禤��@���xH9��g	9tz2ܣ��@v����G%{�,��Ҭ���ق|�Ĺ�(�`-H�uV;��>χ|$�!���3��8`�v���������6%��~��&.����鴀���g"�G���Е���~��/V�DD���)/h�\����oUp%R�Q܆���)h������# �*O��hg�);	`%xpg˯��/k@@���a�Nۤ"i�8B�<ڢ٤ b��ۿ������&�U�Y�&�4ʀ���	_�@�U�)��<�W��͛������Y��8�u����X����w?�:��X~K�cT�F|�b�Z,J�O��))���j���e�j�;;�;��j���Ǳk��"������l������1���Ͽ����Άǧ*+xg��A�g� %8͢n�B��%�:�NIҮ�2�������=��nu�;y�\4NZ1�����;��b��>�f�5>fH_1� ]�	A<2>wѐš3:�T�1�A(P��rh��j���ɣoU$+�IN�Ř^/K�i�����]�:�l�׀X�(hs���YW��) 1�(f�v+��Lb�@G7�ޠ:�-�f��KtՒ�Pײ��s�V6V;�� �Z�&#K�ۨ��Æu���]t,Zr�ns�\���<9O�`IaMr�h^��L��+;�X���K����Ã��қ��v㖬z�,}�c�i�T0 ͙�fch���%����>��R��` }�O�F�e���sV�C/��}����n�s'��R��[j� �T�I�=S"��� �$2B�LJ+�%q����"�F���̘�P��A�7�p������ɑ��L@��'"�l]'��pY)8���.�"��g@o�t�HJ�8�GS���e���%LHh�M��,����k�W���s���)���@<�hݨ�� ��E���s��+��'o�˟�>�:z�~������Z�{j+6	�d�����n��2.�k@���%���$Q{�ߺ����3rEVu~��x�掂����D�'�Td�R�do����2�
b���1E�H�w�|tu��ij�_ �վ�N��<� �Ǧ@K�:kp�k�r6U��K�xz���I�F�-����;�F�2����U�Y�w��Y7:xQ<�lE�l?���1~X���D_��6@np2��V=��0K�7W�	Rx�ְ\�
��Y���FJ⭯���}6(�n_ޭp�&��6b��7��I�ֶ`��& YV��{�Oty���UfӨz߹�����
n:�n�@��2j�f`��#׻�#q&L�{��`펮�&��@:n����c C�NÜ+�QM�6��oQ��$^��xB
��9 �h�Ԅ{�@֭=���ȇ�p�H���!p����l	X|
����61��Gi�ܗ��V,��񐶺.���hCd��qyy�wj�o
v��L*�w���̠x$�����N�}��#�#��Z/�su�?�B���%��;���u��,H#��=í�q>E��G�E/��a��Z�l"��q��.�F��Q�y>z�t!J�������K�^�͋�^��~�\cP�&bU��8��ٚ�>��i!i�Yv܄�$ �kړ�<f�'����~� Rd�J��+]����Se�lT��b@�(�!��ּ��bT�X"��=	<4�-$$k�3{��K>�Q5{�lݏ�M�/8��%��K�����Rw�PH��7�8���;Z�]e�Q_�A�AѾ��K�%�uaQ��6�Vfe������C>�rq�*�h������F 2Tm�\嵏��x�-��NJT��c�"�
ېŔ���/�j�wm�,_ҵ�'���5ub9b)pէ�2��\�$ݘ�r/�Aԫ����`��kw��ڮ��q`��;�)S�,F��Ug&J����.� ��qtM~t�����r�B�h�
��C/P yG�(G�݉2�H��
���䚼�4-�m+ V���̨�e��Ri�;Ke�����J���\���jX�K��dHe]��7�?��$��?�����B4�{��k�7���a[�MIš4c.Heĵz�ēcR�ͯF���q�DփϾ�tʩ�7�/�0�{�T��f?�	��Cdv�.NS�� ��iA3�7��%YI���7�ej��M���Ȣ)'���l�j�g//��ǈ7�s���j��ca�UĀ�s�!��l2�$���02]Z+H���ϐ���������e;���Td�L��5ղ^d��[+�mt���|r�7N��Ɂ8�� �.'k?Pr��Į�@�)� |ŝy�X��U~�kUn�<�U�ZU��&	qe��oe5�DJ��(��>��оV�H����M� >Jt�%Q�d��/:P0���Q�'���̀?�ec�PϢ���CFN����Z�r�/GY��Zv���#����\-�#���h�o�[�n�ΊB����2R��g^�e��Y�啈(ex!;�%���Lƚ7�i�Jϖ劈B��p*մ���I�+k�1��,N6��n�\���&.	A��XE3z�5q�)[�#,��A�OG�[����5�%Ӳ��6~{f��H�f��A�<:�+7���v�/��iWpl�ݹ��
r�32��Ԭ�H�
�c�N9[;�5����ɍ�r�L1go}�:����P�}:�Gg2AގHD�Q&J<� ����!l�L��c����R�(D8�m�@�S+\��z�����iNu�:D�."�᥊*|ר�H�9�{B=ϖ�� �J�6�c+�4RgB~��ѕ�Qdm�](L����V�X�{,*XCa�7�;�z���y*����b�=y��c�~/}~D���I�=#?�$n����[B:d���oIY�೔7Jm��2	s��WD����GcB�\m�l1$�4��u��i!(�����fiĝ����c�����!�?�4]1�lS��o���&e`U�O��׋��}��?.8�
�f'��CP�+6S��nS��	�d�?�B������d޻*,����E7�$�ͷ�-��^���ם�m#֟��"���?VjO�*�}T��݅�4�b}�v�T��D���&�6ȑ9\�X�͗���	������#���0��Ӊ.��5�0��U��i� 5��(�]��j��X���T	��iG��-�{�'�`a�_��-{ �y��8�r5c�����{XS���|N�,K��/ɍ�6�zw��s���S�p�}=Z�֖/����UU�_�&_�ͣ�"n�G���ִ�[�/�w�g�Hq�o4t��	����Y���wnJ,�Om�d�����ز�����$��A���(�QЬO͟.ܤ�� �=A��|���� ����ٕ�0Ԝ]�Kv{�
}�3[�2�|��x��Zט��tV*���Ks�1E&����K��ố{�˳wu&4��L�M>�&�O��>RF�E���q�*���t��&�v��# �ƿ���,L�(�|��鼌�욞�+��l�� ��]h�kƁ*x��9]R�'1u��\��o�@m���hf���mJU��E���L)�q�vM��}?e8�ő���)���`kݥ��*�p���\>�f`9{Wl<de��@�j�8p�(>��;��AֺA!�m�`�����T���p�T)�e���3���>��W�vB}w$;B�Ha��c=k����	]V�` $�+����|n�6};�똆 ,3=2%��f�:�#�����b�&�N`X[xNi�`�Z���~>6�7ld���}�e�����r�z	��^�,;��U��8N (��AIVS�V�Q,F%��2ój ��6IŃ '�u�����ϗ��4�Z�R�ng��iz���o���̦��8|��_io�X�?����389�"�JVA���_�,��[~_�69G��{�]��&Ϙ���S��z@ŀ6Z����e�Ɍ���)Ջ��.U@>� ��B�%k9�V�a\TaٵvX���c���`]R�m ���9m;o��z�!LC�6��¹��ܲ�����o�|�G4W�N<��MK7��G�k����$׵��|�X�<\Y�/��"vA?G�^&�DI���-�Ɲڹ��x�f!�`�������U{��:����Y���ݎ�z����К567 �w{
�Z��ͷ���Yؐ	�������G{&�}O�8�mn����y��%�����̸IX��L'T�D��Me̟/�P�XM"��X������yDk~"�$�$��2����d&��jȚ�(�?�S=�6��r[6�/�y}i'>	��W%�96�Ap�k��`|`寍hg��R�R�b́�TKߔ�HU��^�?/#4��h�yڟ�s��zY-��sk4�U�U��	ߞ�2�5�8��ґNd�V����/�����[��
������x@��f��0Y����Ɍ�7EbI#�j�Eߘ�E��9x���P,���&Ӝy"���< �fЉq��LL�L����gS�����	��v׵c��"���ɕ�I��p���$Y�4�8�잘���	�c�%d����Y�����_�Q�+0"I$�6w��KHy�A�{��$V�LV�iؾ|0q'��P�0����]��1;r'(��u����V�x�H�q�-I'c;���|��R��C¨O�""�ǀ8s*��s�Ĩ��ԟFٗ�>qbt�!V�&��tm�f3Y��&Gp�A��������=�9m��_1��Q�+���m�@g;���Zԯ�4�%�����=�J^����7�N{d�D�p�����#�$�����}c-^bE��PG32������.��!d|΅��hL	T��HE���t��yc�+�*-� 5�#u���P�����i��ZI�:(a���ַr�Ac��$YR�c��$�Ib�QG��z��y7��%�΂�\ee�b���o2�r�D�c8�/a��)
̀D���[��L;q����>E�k�j9Zg�DĂ`@f7�"�`8q��sδUTI|Vp��RcC�#־�k����o�-`�^��dP�ut��2�w;1L L<�iPI��R3lL!M��UC��&_� W5����3�M{/C��_Y�a��A;�M��
��PEu�q\�Hk��������E�����p�$~��&V��%&i��f �ք՞��W��6��D�Q�X{A}�" �׺ѡz̰'�F���Dn�c?�����6�˞v�Ȏ��|I�FǛW#�\х� ��:��w�WD�?ĩs) �-��>����/�ۨ=:�Ã��À��
\��X�|&J�Q�b#\��kQ������c�~���Hu�}�1{z#��ƦGx�����f����#�2��H�G�"_&>����*nɶ���@�0w-	�P\��a������GcZ��B�Vn7���bEg�K�t�W%���щ@%\�> ��@�>��9�$�oXk�K���}�R�V�,�������xv�L�<$�1g���@逈���V8�Y�x%w�A��}0�oq��d����N�&�l��|����h���B ���q���ʍ��/$J����B�qM5IF�PM뭺<���q��I����{�*-�©oxe�U��@V�gO+u#L��<�zg�M�9�m��.��I��r��r��s�:P�]��.� #��X��DU��P�w��sQ������(b�;�D/���iD�C_W���!�XI�b4�M�\qMr���߲�HG����8���6[�6��}!˻ s3VSq/�mHeǄ"
!�a7�m�'y���\�뽐�U�{�ģ�-�f�t��$QU^A_ �߸�#D'N��y����im��LA��-�Y�Lf�?��Q�E=��B����������R����{fL�)��P�'��Zs�|C�s�$Z�ed0ӄi9��T���چ�X��5(h4�熸�%�5�	@h����\	�Ƈs�%�`��D���s��R���l%��l�TZ��;3�Gh��������\���C�c�}|kB�y��l=�Gw�%=��H�����_O�I��O����Ȼ��' �t�gA2��ˋ��H/�y��/�<
9?
��{!� �y���q�)��0�C�pi�]��὿��'���퀁�A�k*��<���h
bĆ"��zB��q˝g���c�<<�?�#�����wKB�*�G~�!8t3�T>v���5˔
���5ԑK���igt>�_8�Ϧ6�����3Q;�dg��O�%�<�~�R�1�}�^-ӿUl��Q�^�r��'���M��ɱ���[\�|W��P�'m�U�����Eߎ�$�XR�*���r��>@�lY��&�� k�'¶����CN��H.+)\v!�w��z$z=��Y�����Zo_+n+�>+��8.&vlOZ^��i3ġ)Z���6zRk�ӻ �z�G��9��w6l��t|%a9j1�'<�<�q6�x����J��C��}�zԺo��`�R�����e���Y�l�I�Z�!A�4���!��ۿ0ڄ�w%��<X7Lp�D��$G�p�*vY���>*���Ag��d&�o�ēZ٨P�� � ,�z�B�����Y�Nn,0�у[��v��´Z2H�׌�*0�rpW�4�����b���(�����3r\�C	x�"�y�������J�H�ʹ�a���ڸ�Z��f������9$J>�-���CfC�Chϡ�
�8��2Pq�Vc\�3��aKZ��9h�����y\��y��/(�z�Qh14���O�>�Z����-��QU}?�I�ϧ_i��_5���p���|EK���ϭ�)a<����A!�~�V�d+�n��Lف;g�q'Լ���;�c0D��; *FI�^*ON`�7u���G<7ʰt;g��PQ͚FV����٨�N�����$%:����
8'~n��vJ5���6J��N�$ q���o�0���NDU�� ��a��ξ�lk�Z ]��G���L�M�!�"(뭃����-��h�j~�Ƌ���n��#1��f�B&��T���W����8�y@Ө�P�>�V�O�%���Q����(̱��(���8���jTGm��1�S�5��3�b*�߃k=?�/�+?D�#�'������|.����,��3gA+�:����F����-��S<��Z�5��b�U������ѤPA�t�_�����0s#�j,�;R1 ��Ws2�7��'1����4ݭ{Ad.ı�u+�*�m� �{��� tr �������Vj&���q�t'���|^j�@�Ìj����em��7y*P`�p�M���#�x���P�W���3%�_R���4v��"����;�e��������^�E�3GK��íbC}J|�AJ!�]Atj��Q2�E1vg�oD��6=�PD7@��B �i��qr�|�R�\��~ҩГR�c4���o	�N�g9hٻ�+K��*�ON�J�Y�P�lp�AwҨ�z�'�ޕ`���/�9���/V�4�x<{i����Qg�{OWS�w"�]�EOË���|�a�ā�4�|� �$��ߤ9Qێ꺫R7��=9����;���3���]��Ln>~�/Sy���jҼl�O�8�a����V���t��{�u��:�T� IKT벇57c�K؄�ct%�/�0v��ǔ���<�����u
�������7BQD3�k��d��E�J��+97�=]��>���þ®A�z��)�����ݡ�X#䘓���4����bI�i̟�ω�X
���BHm��֙����\G_��hst,:��n"kp%`���B�|�L�A;�T�@���[����XqFEKcJ�ˤ-P���A�h"��f��Z�䧶��o=ew��k����ɁG~��)� >���Z
1C���fP,�{2�5>� ��b��d��G���S��UHP4V5� ��u-h�ը��.�@��%(U�Ⱥ��T���D�J8)���2}_�<F�D-�g�fO�r f��]O��o��� �^��/�P`�s�8�4�1s$W�#K��<��q��4R5��Zԯ��f8Q#��z��L�]xE���=�����c��6�C0P�#F��d�+[�#B���&�~�P;�DP}x@����V���1���o�ǹ��`����s �CmQj�z8����A�4���T7c~ޙ�c8E���^nS�WKݐ���y��,R�0���4�h�%+�����e��Ġr��0��5��l����U�)+̴5^�;���0wI��; t��4Su"A�}�_��E|N�>(X֨�J�Ԃ���r���{�Ń�L�1�W\mF$�?
	 �*ix�R�6�1@�. W���2>ג�6�����Y�1cb�:�V�l�P8��u��rr���}�M���sP)�H�_���\��g�����S����P$�g�:���#9�v���h�Հ�B|���q6�KJs>�5�6��}���d���Zǲ�O����[�.����t�ߏ%LZu�c�Q�vxw)�5c'$|�u�V����
_��k���:;�q�W]|�xX���خ)���y�}Q�1#�)����i��"��m�B��h�ʩ�|j�dG�%�+z ?ߵ�k0�%�[���Μ�k&IO[�G�ﺠ�2��o^|1�hNq�U1=��;�(�A�qE��+l���׮�Rn��į�:!܈�P�||�>wS.�^��F�J^�)�OE��V����I�m@���	�5�6�m�u�ȶUT&ʫ��7�ۘ���|�M.�)eY����|�=;Y�q��5��4��s��5��16�OAz����	a����M�X{�1�۝'�D�B�E�ڪIY�n5�6�h��&�|�y�(cO@�,�9A�A}j�����ѷ"Ӂ�3��~����A�m�ʎѨ,[bH��"F�8Ϗ�}̨�=���ÀCڄQY���-%i]���s�57)�ϩJ��E���#�K�|�L:i�S��'��6h&�^��"�iS��ˤ�.*�|r(>�]k�-�c�w��O����dZx-;�$���	�ނ��ߔ���C
�qf��&���U5���2�hB/�w�c ���Qbt�7'��ɥ��y/I�}]��3Z!���aĴ�`�=z>�m�~���Xx����ÿdyy��+?���i
��#�Q���m�F��������V	���+N��c����&% �|�����c�z�wva�X*��#(*j}�0�/�t�[�JFB3��ӳ�2$���`�S���J|��{	�~�Y��=����?�����\[Q�͒����Ƚ��� ��S�	A�a���\5�4�-b���a�Ā|-�����uW�������3�"H�iE���e~H�����h]�s�v[+�.lfF
I��ի|�����^���+2����K��&ߥ��EU1_δ�M~�v���ف�_eiav�.]1��$����tn<�m-׻�M�_i࿫F����k��k���$�H��.�#�Y���Y�.0wlFX�}>�PQ���������n)�焥��ӫ�Lk�*C�eO��\�U��:i/�x�>O�� /N��co�]��S���P4R��c$��j�/#Ѝ'��μZ�Q�� P�YL���ҒC@�1u(�t��o�H{RI�jl�����J�����,�M|�2�����mi�% ގb��׿���
~2��ȴ�c�� {9�|TU��� ��-f�w�>�4>-x���a`+���ƭ�ʒo������u���ۛ�w��߰��^<�Z��s���Ve]�ƭ.��ѡVWVi��w� ���b]�|�g��~�o/��tS���!7*���	W�b	�ܡ��LN�DҟW�[[a&J��;�=��^٨C(��5g~�-�˽�k'�(�M`ޝ��`ro-ÿ�<l3+漹�����bz���
�9o��I�J�Ġ���A��M�|,|����Bv�Y�Z|��Tt�m,#!�:�KqA��ڄOE������OsX� .��IN}x�7x�'�}�˜�fٞ�H��/濮�RJ�%�ܡ�V��,v���V�q�|��Ǣ��9}H_����RI�P,HN��f��$xz��b�>c� �9�A����*4P�����^f8P�=Α�mA�m|t�ő�Fw���������K�����X�� ���H�	�b���wLmIW!'o!1kh{���\���ő�FeW^�G��F��{ܥ��}�Y,��lSȎ�	'6��)I���c,v��&�Ǯ��_���]ޟ���?���
Fn���*�s�I��QC���Z��`�@��('�{�P�4�\~��O�����~
 �CA�O��~0<�h{����;��H��N�"H��;��j�}��GZ���A�^z9ũ�P5��E�H#e�x<̈́����kg[�b��[�-⽭P���[#l���TO����V�����S��;$�@]�&�y�Q�;{V�����9��_���	nXi��?�+f�ɝDn��8\;+)��A��Z�|ctJ�i��3HE*�X��:LO[)o�����zIh�_��i1(����w5BC5�M`�tݪ�=D�7S(;��HP�W� �R��^	�յyZ���^L%�>F7�*�O�.D3�~�������o�����G8�hyGo����:�o��ѡ����XNf��P��v�&�����C�M�e�z���x�"�l��!o{���M<�{ݥ9[�*~1����	�D�Z�W��W| oDҡ$p՛'S_����a�HQ{��Ù=(n҄�8������#;Ib�XlxVHYEB    590c     f20���^0DZypW���Wݣ%��$�trD��!Z��w3�l,�f�L�b����g検�x���<�x���`�bb�۾4Ԗw��:q�%����x��O~�\'t��~� "��F��f����>\DITL�P�\�e�@��ˤ���]�[P�C��BD���|�B��.F�eyB���'/�*˪���pSWSW��MS���zOAGJ!rZm�6�	 ���x�Y9�`	K~�!
H�2}A�>oj��+���ٸ����/P.Ƿ�Y
�긝��bkI#e�D�`J��p��l�mJ�M�V���x5�9bp}-�oTU>����>{_UT�%�s�fd)V&�g��Y7o���[�̽w�o��	�C��^�x��:vXl��4�y�{Ƽ��6{B�@z�-�I�B�9F�������p��������M�}�(��	�����e�i�H����=�c���뒩dѬ�E=���բ�-}_Y��^�]hA9r�˲+ R*6i�X�O��{ Ѫ���6�� �s40昳���PSXj]�\}6�Ysl�f��������sT�lq��ٞ#�8���KR��qw�k~��q!�^�uE�ZO�=�BHnh�
,�Ȭ�w� 7���W������r�C��&(?�1�C'驡nzҁ�6:Dtw�K�������\Q�t}��3�u4�'g8)�Q
�nC�C�ج4����Esm��U-�%�G�9�t�x���,�v���RG|��W�d�j�����.y�cd�Ƒr5�M��>M�r��t��+5�V�t�{��'�҈n�]j�1���+��� t�1�.���@-]D1 �^ (���iLKpI7G��w��B�69v����XHf"E<:d�i0 ��8��$q%�c�>�@v '#8��+���p�����k�b&I�)24�ai=�LI�)�B,	����A��8�.'aA��ZV�r����h�8���j�&p1�m�3��p4z�2� ���$���v��!>�)�h��m>Q! ������$�7�c	E����<�k��j5�.�X��[(HtXW_�Є!��̞J0FU��o�ӄе=ԖFY�0�u8!��x��-�����H�f����z�x���+q��N��R=.+)��e�CO��\6�U<w�P=ʘD ��pl�v�ަ$�68�=X.�>�Q�h0E�>�C0H[�[���Hj�-�3�����HtU벱�;3�ߡ��r�'�1�wq�ګ�lx!8v�us��.z�G�`��b����#�T����4s2�������JI"0mѰQ!m�����q��A)`_��*������� '�x��!�ԣIk������FE�[[']����MJ��k���=��).�u���![:DO��*�^{�ǳ�I����fR��dG���'΅�����A]���B����;D��d�c����/x��`<w̽\���M��/L�n�Fs&�L=�I�}�Gp���:���?B���Bf(o�*	l�o�͘���-�m�:@ZT�\���#���e'ʹԴz{J�(�?L��c2�Mǌ���l�*�yvA�����z�w�~���Y0���{�A�A�օ+|tuQV�!a�������!`�$����ъ�P��Ҍ2��2��%��½��o;�=�y7�e�"2�ۃ��[�A|��_�m��>Y�R*��@Zm��.��@:��|m�[l��&�L�G�^�+�P�Oɤ�4�}H�%"��(�d/,���:6�]���n���U�^�&P�}C� �X�@{����M�c4��P�F�L�^�)�:�Jv94�i�K�i�؃)2F:j]Р���D��ݲ"��dk�a�$\g�o�V9�y;��
\7��6�>�$7�Sr8�ܢ7�s(n�� ���Ql��[�nD�T�E0 �c��%ę�s�ۋufs�eon�6��f���FR��y��� �7���ƝsGE\����p���C#����,^6���uq���f��E/S�%�+�BOyΰ?�V�(��0�`؟"5ܓ$�F,țW�$.Ҫj+�b'�~���؅�㷷k�O�v[D4"��;�����y8k��ݨ:� c3����OȶΏg���d&@��|{�$ ��!��eܪDL]��pFGY��e�Ĺѣj�u��vy�D����s�9H �+\Ed�4#�=����QIVy��B�ޞ�b�]��%��<b�˚_��6۴� �[�3�o�W ��h��"u�����Bו+��:��Q&�11~afB�����S�0���	�ln��_j��b����:#5*��kh%�|?����(cos���dnn��T�8���"m�T�f�����ƅV9��7{P���3*�-$@�7� ���:���M��+b�?��`m��Ѹ������兲����T`���j1�+n�z"�iM@�l�5��ix����z�R>^��L��Σ��[�;���D�J�#y���6���``K��I��y�����ۀ��M�5R���U*�[�eiW��W�8Ӏ,��&�y��,��[.T�*I�hK�yW&�8NdS�_l��6Y+���N�ގ��B�[q
�2��AI/�@᭑cm(l�H�tK�w�v��ɗB��Qr�y�x^��@� �o�"!.�n	{�v��%���fn�6�ũO6�v�C�0�Hǎ��X�RסcC͜.c~������D-�����S8�
�>G����Cv{��PC9�:��$`�O0��_�<MeW�ԹH'p�$鳻"�i#�h�(�z��'\x��E(������.�{9��R�,�'�
��>�F��Ϲ�%2}(ꔸ���G�L���^��ѝe��N�vu=��xB�cݤr˳d�~�NRߓ�!��42z	�c9���p9�Ov~��o@���u2��J����4�P�og仧(����_����ZEȼݽ�:d����!�<��2�������֮~ �e��f���,�}CXq�,���޿�!rc���q''9oA������z@���E���fR�i���0�;�O��$��0=� ��I�1S(^�K����6�~L��*P�ёr�}�0§�|�L` ��y��[BV�aU��[�Cںqc�E��A���QV�\kk̨)��DY�����H�=�GQFrK�@�����"�Ow���T��Fӧ2��z��N��G�u�ݰ�vʠ5��s
C��2d�H�?e��s"kQ^d`�Ƽ��3k�[��3\Z��y�����mYE�Dh��yl׷��+����M���Y�T����9�$9Z�'r ��eLA��zk*$��&��`'��9ĝ��o�C� Ԭ,zС<O�]Cǫʨ��g�1��%�0��b��;d�|��<W�C���(����M~;�[�[f�j`N����y���w�����5�i��T����]��pP䳭qr(��P�O��c�w�Z�U^�ݭ�H=ǩ[�O��Ѣ�������wd}׽�9��	����&�h���Rn���$�E���f���%��p��K�^!a0Wmn�@��}r��я�8@=w�'�Z�]� ��b����Ès�em�WLݞE���)����>�>���%E"��6���Q��v��8��͝������;�zQ���v���asK��<�QP�/�KQ���b�K�K�#Ҡ{��ɭ�T{v�i6i��JbA���-��-�F�⿃/�t����ڟ ����/]]��v,��|�|��g�q���`�3Z8Ҹ���A}����7��䓅��2��,��\�c��/�>�F@
����=��J�x0�d�Q}Nn�\C�b��]��H�������_�Y�O�%��=�܋����