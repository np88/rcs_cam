XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����ek��#@�&9?6(����g[��i�lM�{�PG��I�3@\���gn��{��/ P%�m�b%@_CiG�G����?�H.����o��8����
d��3�5�|ܩ��	�B>��d�f���^�����r�.�C��\��A��>7lr}	��lZ[�]��0�R=�w�4 �:\��#Y����H3e�I��pp
*��t<��%�L��N�B��oC	pp��K�G����pW~�ėy┉�v�Y�9@��������k��\h�w@��îf D	�e���\�|y�k���L�￦�-H$����F�;�	Y��]�+Ɲ�3#!rX<�w�������;  �p�c���>­+u�%}��ʲ�ʀGV]?M.-{��K�5��M˴u�W[X�L���N�6τq}�E�K�nN/�|i���pՂZ�n{۾ZC�
�Q���_��s�ܝ��_����E#v�6=W3B�Mf�2�]�Dd���)r`mφď���/%�	�����~�����]����~�X����ǚ:����`,NEa��K4�U�O")�!�1�h�g�� ��=Y�����0�J��Ā�m� 	)9<ՔCu�ͅ|^ވ���4�h|�O`[�<�0t2���ݣ��	JZ?|X#�ug"�q��-�޽*�>+9R1x@͈�q�C�(��!�����xtt��@k��B�%���9�B٩���T&�x����R肅��Bp��iXlxVHYEB    fa00    1950�3��qtJ��:}�ܾ�>!;�u�b	��e�3T�>����J��Y6[���d6Z���N:,,����DKT���I�s["XR�9T��ij4����a�{���
�A���~����V��ҡ��i��	����xvҹ���y�[�����ȵ�/�P�y���4�0҃�e���H<Bjd[��}:��E����'����ſ�V�ɋa�q��.�I���B<9?4��[;����mj��=�k|#v*�8]���#h������b�}�|h��%��/^��!��W��[��2�Y��8_���#�s����vѦ���\�v��=�V.��r�rfX��7���uz3�ן�F��ܒ�N=���$%�6/�H�2�;��h�^���w'v�v����`Q�o�m+��O8��̳�`B�NX#3�y�(�Ҡ�UK�v?���b;�V��7ݯz���u%�V�i�3�,�4ܽh�w�$�կ�g����L��b���Ǧ�������e��H~�n�]��Z�|CΝ�YW�{|�Fׇ딲�G�#�;�<�O�mۜMJ���!z��h��3�%= haF���Aó$�\T��Q{�⸪�45���9L��TN�l���
���_ʈs:K;_�3�zy#�ԝ���H�����f��BmQt��"�MQ9�G�E371�1B� ���)�Lq�����q��A�4$��u$_�u:q�-
m�?Ͻ�n��^��A�Ƈ��5�ٗ�s�g0�#¢��~�X��Zʔ���͟d���`�FȈJuu��B"����n�Iȼ%���T�Z1%8N��?Uk7�%fL��F��g�_��h����s%:�y���#j�P�����:|�h��R�Ss�a�� �"� ˘��B�\�7^��R��ռ;���&(��s=֪Q�g�bZǌ���t���4k�@�[�z@@nͣ)
�W�a�AK�y�:�/\y���g����L������TfT��͹����%�	8���	g��_�ʳ�o��i��k�d��>2��,��.}�A�w�-{�̉�y<�1�9Hy/��g�ĞAr����y4 �[�]���A�O⽂%�|g�W%rd;y8�����n����mz�e��	��ٙ���-�G���$/7��T�4q25�3���6(X����Jm)ƀ��h	�̪��дL`��A��H6�Y�J��;q�H*�1~n?L*k(�s[�&-"��H��Eğ��u��f��y�k�z��>&��oF2.�Z����H��ϕ�c���A��`,��}���fP�e�q��}������KS$lI��^��g6���l�'���m/�[~�O�1Ǒ���"�m&d���8}�4���O~�����vw��9Ɛ���J��~���ͤ�)d�p�Po��rDB�ZPN?�~���� {Y�&���9׍���a�ƫ/0b;��y7p<*(lK�Oq>T1�Y��v��5�C�����aeԇC�b���<���C%�4�Q��,�-x�v��8Ou'��6�lZ._�]�Q�S"�/\v~��6��d�8oX��P�Bcd|��̼�9|��~x�Fo�ơ����)gThm�Cv����։C �����ǹ{��E���f�Dz:˅�v�n'���T�vV��c�%SS�^��~�Hez%<{F����A�sV8=Ril]^�`�X���*���&R��`�xS�<|%e�*�?b�b��)��q uX�zڤ��/Bń�L%l1$���zmM�a@��^;�~j�K#W�R�?�&�B��7E�:P���ZJք�8j�>�M��d!IVc��D���*���lwDCA�l�R$P�{{}�-��Y�>��O���Nq�ИX�3�e�B�P�USf�lo�xW.�A���r�m3ueٔu@��V
f3�dM� [�C|���-a='sH~�֏��+`�4s��v�rO^�L��ZBQbL�S��)��*V��i۠Um��|I`��K�G�� :\5��?�G�r��`��oS�.��X�����(���yd�N��	R���罊��g��a�loc>�U�Z��:������C��b5C�`�I������_�"�ti�/�I�����$do�����Or~&��P*P��wE��t�z��V��p1�s�sqOTu�\V���a���Te�"����@ᖂ/I[�����3��C���6��÷�4�EX"HS���$��Wӳ�@��~~����X�6��B��[d;=�c��8�t��&h��_��"7c��2��E��-�U��U�*|�uWށ�1�>��F�N�`���w�$mS48�G�����)2!sj��&�ת�z�i��A����Q�����;�J���Z�l�GJS�)�����n��4�JRǠP,k	�[A?99�V��S�-IgK5>7h0'W
��R;j��[�B`�����HH�\l���zd��gw�╋d/��ؒ4-��\a��([SN��Eu���1��IR�h��J�i���D�G{�z�.vLΜ�?\1(%u�HF��=a@��C��+��P�&�5��z����N�����6�A �^�t�qGsy�(/m�MgU�ڔR���^�%ܨ'�p)sQ~R~�]D�9�@����%C1���ŪOe�~�yљ�28ۛ�@��ǽ��W��Y����%M����ց�<@q�i�G�H?_w}�{�4��r��߆�L�5�K��B�@�s�v�?����/��uA����-�������.u|���MzA5�nD�}��_6͒h�l7K������`���c�T*���+��X}3>��c��ɂ<����O��ňT�l6߂br�-��^��G��a z>�����Ӟ�*j���j��CZ$�=+���{�W��'�5�5?�5+;��Uy�Py�����
>���/���c�N�<�-8>��xSV	��A��P	a��`�S�c��� O�P�8�Y�kpd�2���M��Ms~�w�5�;�ȶ6t�G	��<�ˋ��jf�H1������I^ʪ�TD�5n���i�mt:��Xx�FK�k"� ��J:�Mc��ٴ6�{�}��g�9����,Z9������6�|-3����ٺ��s2���[GH����vו��J+ܲ���+����*�TM;��Ț�ep��V���ք������b�}�����,��kӈ0��@r����C�³[�/��~[�ω�L ^���}�.���*~:ƋR��c�p��H��%���NS�ڰ����s�l�]�3)/��V�	���� �ry~g\
%A��^��H��j�e�h�\�k�1u��YB��Hs�,�d�[όj��ob��ØW�,�X�柟�WN�vO���U�,��]�@���AS�ILn%锖?K�f���/�g��a<F� 
����I��
�(�0���4	KS����'0��+�HYV��	�S���	b�U�1T=Pۙ��'��YF���������z��s�'VP�pSr)U�6����e̥j�L�����r�@�S�)�˲���V�/`o	��QR��$��[ch$�=��(~&b���k=`N�:1�|����O�F��w޷0�Q4%V���q����j��6H�NŠX����Q���
�I/M'��m�M��/����]�[����sЮI��ǀp������e��R�Fn䦁�j�E�m? ���|��;���
8&n�Q�d���?�Wl�Wn}\�ޥ.o�C�6S��<��̲��~�?�x�����s��m�fB)���W����nE��w| O7儩��Q+��7#���e<Ub҄F��p&����0�oV�,c�{�&�<!�U��~>�\�7���KDq!�yM�h$&A�b�z9c�Z�TMz�i�?�;��l�'b�����@���>�1�p�m	O�<��W�2����Sv�%Ns��j6�*g5�D��<�M�A,�f���q�{^�
��&O�r����p��)��ę�,�t�`�[Ѡ�80��}жP8��?P�/�K�u�g�n{δ'��4D����Z嶅��궉�(���̗���A����d-�	������U��L�m&�=hS�uܧh
7-/���Ԧ$~�l3�G�fh�)t��Y� �V��@Pu��o���0O��cI�)ڿ�zR�$@k��:���S��D�2�(#��a#|ӿ�kmz�W��W�:ϭi�{�z�̓t���,�𒦙�Ԁ,�S�t)(ػ��̠ �� z}�c���t[E�b�O����g�=|U.��ә��A�c��ᥣQ]�5��>:��8-�ƺ�q��f�2P>-x[s�[�ɎLp��;ҩ24��~������d�X��ϸ��9|Ǝ�7��WdD>��s�nw�:�V��fL�p�M�Q��꺜�!`�R�Dy��(�fP��v�<?��}4c?u���Z�tY�p�<>J.��3W�d����=+T���P���r.9��yp7#��8�|�}U`�G�mcNS{K���2�� DD��k���>�`����/ѿ4MQ�&_�2��OY��Siٞ�����{���5g�܉�V����C*�ҧ��;{\&9�j��*���՛�+P�fX8��B�a6	,K��~����փ�A�*��;ЗRC,.艰H���R��z�[��U��w�O���N�|\ﶿ�XI4�^)�|[���*�˴X���x!!܇���-vfJ��`xy�f�<��8�	������M7����\rB|r*�%���V�|}0q�㘢}n�Ow1T�B���������]13�!^Ʌh�PM�L�4e�i��k�P~�x]r����u��?Ӊ����$=6��e-s�<}u骰"��c���%$� *:�c�ڰ3�_`C���G����c�=���K���'��,��W� =&���YAus� 0L{e评�A1���~�Al�����z��Af����X%�F�?Rͽ"N�,�{2Y��4x��KǛ9͢%cw�E�yr�� `%W�o�T �/Hc���SQI��D � � �j�5K����o�ҋ��_�w�� ���Ni�Z�bNMd�Z.�AJ(8�627�0���|����UO�!����+_��:�ٱ��!d�4^���S�������46Pz�%� P=��F���{Ro�$���>�"�:k�4AEJ��9������)�2� TM4@�g��Q՜��x!�﫱�	
䉅� x֋B�:Mטuۊh?I�0��C��s�-��}eN��8r]�� ���b���7Q����_��ʩtab����F�V����YR%J�P+E0N'Q"B�Z�����ц�Ƚ��.��{u�I2g�DI����x@,EN�Hb!�����p��5��0��BB����v�L���d�k/��Թ�	I7�*����~�nW�N[�nbᕬ"�0�˕ϴ~���ɯ���{�̦������Ǧ�uL6��1���A'Y�w�M)�-f�=f�O��������R��*�`[��F[P�$+U��k�����'�?^����Z3pM3UB���
ay�v���B�q��l���$؉�s����X���2��%w��NK��>�H�v��j��1�J�_���B$g�3�{����@x�6��9#���w<C�v��x�8\�yq�Ď���Vw��W�A)Z����57gR���#=�>}4G�4�ȗoH)�tkN�o4�;y�Eyޛ�j�������{N�e(���"�����'����7*��ړ�`(� ��JS�8͝7(=�n(,a�e�4�Y��57h��^F�#OY����hI�>֍���8�f���|R�
�' z�+؆�rLSM�q�y���C�:x��w:���4�T:L��?��"?2�1��*/K��2~��S�)D�M]��+Т,�(k!Y���[0���B�����0��"�C���}��!�gKl��V4��f"߇a�_�HTK��~$�r%�,Q��;��5�_�!>�X/^m쯮�U��f�#�&��;z�Ä�(an4��	]�cy	bH��-`�����f�64i �
b������s�O>}�Ȅ'w_Wp�����C�i���6��`�����]ǔ��g��k���4�[I׷��<����Rs�o{2���a$�p�y���xU	�����+�FTI��\"�Y�8bX�5�l��0d��A!�B{�Y��ma�w*��'U��kA��n�|����%�H�4f3���K��;�V3o^!I����s~�x{�����x���`��|$���*/Q��W��${-�c�_�.0'������j�U�sȽq�+���/J��/��-���s�Nhq�a�d�7�����-���u�N���ʘ~��i:(N5)�@C~��c�r��L��^5�).h� Ҥ�k��*܀��E��f2�ږ�[+��sƞ�$XlxVHYEB    fa00     700rCѶ�����#5��D�f�%BN���ڋ�dl�/��(o�!\�Q+-i�H��:Þ��2�.�l�Zѩ�fO3�~^�����췯�O:������A�sa}�����]�zs����2�LO�,n3�.�1h��!�p*�r�{p�1���wJZ�[���+���2z�>�~�CLMr1�T
"KY��A�o�Y^Z�ih��@���y��Vnc>&�A�@")S���sE��x�b@R��|B������(�v��7x6
f�3���;�=�xc��DJ�+4�gW�������8�9�m�Eܔo�ĘH@��h7�"�%�g���.ȃG���;b3�R=x�$D�O
�W�}�)^^���������U��sh����d{E� �;:�v9�U>I���~��\�h]|W&�",_�4 ��R��h�-Ӛ=H������;D��:#���Dn��YVX+��Qx�1�����b��V��h��_ U��p^PK�&s�]Ê{z�GO���xq�K��'��!�$5W����t&:,ȑ�@����!�j�vn����ڛ#Lˇ�49��H᧰������UԀT7�C��w�u��t�_]BAv,�/������M���b��yg9]<`�~�T�w���F����:��kR%$֪��$0J>'�G�!�M׈r�7�w��c[���1M�'��G�����Z����'�5�)W��N�Ze�sfd �%>k\�;��1��~�Du�e�L�h�N�_�Nx|?��������>$w�M��,��;Y9Hԗ[O����rD�Wиk�_���Y����Uf+�}���Z&�3zf�&�Cܢ�<��L��B�{psjra׾l�7�]�*���+��=n9��d@��Zu�΃L>�������K�*DXIt���)J��������D𖣌�f�CoB�5bN|�iUb4�t	[yE�%�H|P�$Q&��@I9	���|��.K<2�l"܈/�$8}3~'���}�-�.�/����8�/���-ӝ=�ԉ�y�{Lꦄ�2����(�N���ClEI���V]�͋a�zy
eWy�R�k�F�3�0�-����k�=�P	�K���8�)��d�p�L}^5)�I'��t�e]�BY������znz��5��'��D�%8�����~i���||�!�D�t�!�z��h�tTn�cg��L�n��t��o�I��-q�q���Lyzw	t*X��R	��7[k�������:�Z���D�"���C�R���P�/�9�x�>M$+x� [vP�`�q���p'$�}��4g�4���uo8��t�g��!kD
���?�X���E\C�ʂ�����H<��� P�
u���hpKK����.���V���4�vwn��g���9�G^I����몮ݼ[�Kl��p0�ȋ��Y���;g%٤.��:/l-�s&�1X�yIw업,�x��ns�K�0�_�,�����ꃦĬk�y�D�!�3�/U�,͞����4��g�!�'rO���c
���9�:a�Oҷp���w�Qi�{���#��T��s��|�v�|�����j�����j�ӄ�8E��G�[��E�G�{�R��R�h	�����7h����߿/N�W��Tz,�Zŀ���a��M]I�r�έx��-�P`�%*��������Xf��(:]#�(��=���'p<����Wi��ix���)ӹW_�l�,�m� ��û��F�F3�UǶ�#XlxVHYEB    77da     a60���5�N\ǠN)�js�����J.�"o���eU��KEUk�X�ڃ=L<g�Ȱ띻��\�<�K3���-�E�A�(��TC�c�1���5b������j+�i�9��k�B2xQD! ����.r��%�,���3�Y`}sx��&9� ���d�SU�I��S�aX��wp�ٛ���a��{T~.����a+f�O�巖�X�	v�i ҋl�7z��mHD�0��C��%�7�C��b���/��<�>�U�Sq������?6O;>0��x��j�h�	��OpTQ�߿_~˅G�F��Y�*�HG{��] h̙��2B��3�����UI���=Q@I��3藖H��E�W��y�e���I���><�� ҉���P�y|f	K����r)�W��H�!��P� �"1���8E�i��TO@��ɟ��dӶ����(�H����in���ډ1^4�	�d�|[0��T��՟����g���h����Q�{�&��󑸓�R3*g+}�R�R.hX[��n��z�8���8A �Z��e�n���!���8W���/�����@#�VVB�h�O�����L�0�|�o�1#}�s��Lv��&��e:,I���(�ώ�q�� ��9�������0mo�u��DL��0��X$�so�A�Su���n�Bߺ.�I���Wd�ρ���P�jL|�D���Ze'�{���i����:<�K�����#@��V~&N������)@��??��7�/,��4�`A*O4nuFp,�����oo��K���m��Y��C��o&p�!���a
��c�a���~��5��+^+Q����"�	��CЙ҆6�)�j�\��U��#���v��$+�j���Uu���P��q ���Ɓ���R��^5�G�Qu׍ ��D`�U#���̶��
�l+�+E�-=�%󆸶�������iČ��Fq8���FaIL�0����<���d���y�x���-����S�s����m$����G�H�G���>�/^���"�� g��")�9�=_L>���Es0a2��8{Upgz��L��ވg�X/�G�D�_������o��ֻ	�_��,o[+�&*�>Qߏ���>��k��IX�Z�a=�~���#/�xܰჃ�@ѕ��5|2���J��A�u�i�Fz�J��e�_�\._)��Zg67/�Rm��[�{��q=0 �{̅�蓦�RxN�Z�
^����8�$�|]+.�qMQ5��U��"`�%�õ��ALWm�@٧R.�����*�5�ƽ�.s�?P���Py���}�t-$�t4�O����y1��ղg�,���7����u?�c��ç<��d���ɑϦ��K�ắ���D�s�R��m��M�z�|�k�v���dc8iӅ����f��2�x�n��|�<L���~�ver����i����h ·-����4gu�D����(l���jZ'5-�Wb�͂�v����K�=
�W�˃_wb�y�*���\�w*6����|��N�`��W,{p��n`͎�h>��Y(jE56�������ǲ�����O�h�������S����Ե
���|�j����B�6�Ϩ�va�WR�j�@��%��؀�|�q����f\��@s�&HϠ�U��e���4�����h�[3�M�5+6�f����n����HoR2�$CX�g��i|��������L���M�����X�Qĸ���'&�������+;�i*R�ȥ�u�jd�gt�J��r�:֙��t�"��j��������;?�ͻՙZ�!h�I����T��|\g�����@�y+m�!0Td����Z��6�%EY+�#v�t��1������6e���6BJ�?��V�
�d��A������lPi�^[�+�����D��^�Π#��C:+�?9�5�/U�ޝ�k<9�^PYK<Q���Zm�J�"_���D�
2C5�4����l)~R�B�b�jI;���wf��;o��VG�A_�cbЁ!bM8��K�!'Y����jK�y}�εo��Pt�3���?&��g�U;�¡�˱�v�/�8�*u�g��K+�+,��=��lK���A��{�/�G?Q�%�2��$ׂ�WI��͏t�o���v���Z�Wy��V��cqG�Dz������s�`���4LCK��S�=t*Lk�����+�i_bA)M���o�U#'�Au4��c�f�����rf��v@��@k��Tޙ)&X2�-�OzBc�9��q��-5��,�5BmX�R���׻�������_l'v��Q��q(�Njv�8w�X7~d�����L�L��,x����@��_c|s�tkk���M�,�#���o�~���Ȍ�Ls�h͆v��3^�\b6���9b]�V����@��qў�f'�����G����K�=0 ��~��Ww���P���ήQt��A�JMh����;����S12ߡ�� N���2];P�Y#K���$��@��u}>���O'9�)��zmԦ��M��+@�3ǫ"�Y��p�p���ẕ�_���.�Ϊ;���������s8א�i1c��8y[����U��E_�3!w_��!d�