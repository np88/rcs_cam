XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��@�j16Od�YviX`���g�sبC����Q&#k���"�kr�>d� x��t��4Ӏ�U��ͪ�c��x��Jˌڲ�~i�LW�{��ڦ���Oe�a+B%�"#ދh�2(T��k��f���-g����V�0c��~��B!|��Y�,��t��uoh���]�2+�Z�����d�P���#}�θA�� �}'D[|5�Z�#�`w��A�̦�|`��ZN ��-[�k�J/�5��
�-��(f�� l�lۯ�ѣ�R����ͷ�o+��-�v$;�F���$���T�}m��ƶ�w��d�!��E�b !���u8�-1�n��8�5�����Ws+Q�i�2?0fQ�u������*��a���F����$�����*���#o<��	�G�����bz�a�#J�s�y(�%4�瘚,D)(�VD�j���H R���������y��U0Z������'�U�����̼Z�r�;���EN���Aj�b�]gr�q`2t�,0�,���Cg����q������Q����c|c�7:�"��n���i��ښB)��J�,_ҷʰA�M�=�6܌�]�O�3jr�+��\%/�!���)�^?y]�pa�oL�����{��>�F h.O�X�,z=a��^]eWԺ���Q�����ȸ
����K�Q�U�ׂ�([���Q
{R���PF���38N�A�C��3���o�q<ͳk{⹆�'J�3�P$�%��Z�18��9��)Qcx��8��Kye��D�XlxVHYEB    c3e8    1d20¯�P��D_��k{�x��By>C��%�{��f7�l�^�Ŧ#i�X�/�I���5
v逌����J��}Ǎd¹��s��1�\u��5 �~�0Q��ӮŞ��K>���������;��m4|�=��J��%���)v�XG�|�����<q���ת�mչ�h� s�"t��Ja< 4O�4}��(u��re�,a]/���!���Y�7J�d�XN鵬���"�� o;i/�E澁��5�y�rK�$-���KI��?r�l�<<����SyH%���G �f�]/��C
�G���̀�~���o9�(���uX�o�K��ڂDa�G.��92��ot1�����1>G���mU*x������@��#�jQ�!,N��
=F_��~���Q�Y�h�����9�5�� Ѡ��Fc�
!��:'��j K;�2#$J"`�s��^IN%:�<=���%ob�<+�n`1��3΢o�S!�'�<xc6���I��d�DLӿ�%R�(���:\'<�G��� 9�g��G|�*kc͢@���˶;}� ���H��6�:>O�C7)��ҿL�9cC��(.u�>���?d��6��7{y���b�f�A����|m�j������JX���.a��GA</�h1t�����%�&�܈�2�}W-��2�*>� ���~�lc��z�:� F-�
���^�#x�8
�z��;��2�
i�����eV��2��Z���`r!I�,A)b��5�=z6gɉ���ο�o��W�v�JB9��cCn�(sQJ~�����kw��ZB,�2��|�cȲuQ��{$�|8�O�&z<i�f@�;��Bu�N�.^�D|y3�/GÎ�}g5��[S���(��!�h�����)�D���n�E��TB$>�:�@��\*�����Kx�Q1�h����[����x@��!p��;�ѯ� �s��\�/6%s�0�^_&��!`\9�B��.c_�V܌��a'm�z�$R&���cp���sȨ�}�Jp ��g�����]�$F&�T �_�d�3�U��>�YG�N�X�`\JU¯��V�T2��Ps��#�̃�¢w�z���'��	l��~�	�CK�H��?3Ѽ�El�WߨȖ�O�Fn:��<��ܖFc�1	-��!)�r��K@�o
�8�;���C�o�#���$���[���*b)p�f#E�3B6K�.��Pwܙ��z��,h�k��إX�J�Ӌŀm����@;i�8�M�"���N
�nl�r0�b�������x�3�v;���7���&A�D�n��-�jҮ_cp�=�����d��P���@�s�Q��q�[���T�El��3+Q_#FK�g��k{S���A�@�,��������>��4�����뻕���bmYhJp>�������eW�q���z͒u��Mk�����f��~9���ag���׫���k���RXN�s��7��ِo��D6T��U����Z)`�	��UȐ���Y���@�O"��N��H�3�kq7��bd.�pO����&�'	�~�G�7��C ��ANV`s\��P�Dp���T��|"��Lȋ_��=�!�:�j�����|FX&�k$ZHT��D�SNȲ��X£D�� ?B�e ^(L�l%1F�W�� @�˗S��p_��r"�9���/yM����_^��2Z�B���yB�c�j�t?��<�B8ik�<;.ϨR��_18��sw.'T.%�q��mg.nb6��~y���7K�uY�ò!vˑη$��j"��6��qd%dɌ�k`Q�� �L�^Â�Ӫ�9)�\3��}VC��θǣ�Q/?��jIٿx6��C�!�f5O�@�n���m��U=L�&�?�E�����O�c�x�|�z�K���_ҿΥ.i>s�F�'r�����ϲέ�r0+u4"����;�g��٩6�ʮ/�u1�G����B�I`J;EἏXݕ��q*���}�S��.�Ў �O'��[�E�>�
jU�.ڦ��W�ϴ���6%���!�����\Znno@��,�%�v�YW��g����k����c�Zq��%��	���&6?m��&v�ޗ�#-o�ּVnIB�R�p�3
3 ]6��
2�'E5�#b�~��}���R!4�E�~0%�!>r�I��	���j&��Gج���"�~d�'uס������H�`f3�/�k�=����;�"�y~�yUn����Q��^$�u�h��'�bCZ	�߼�WӋ��D,*@�p����2 ��{�K�E^����y}��E��{�#��v��)�s?X削r� ��҇'N��M
|�?���3�)�)G0�����T�Pʀ�jQ[���OQ��V�'o #��Zq�U��3l�|Vv{Up�p:J��Ռe>o퓺��i��9μ���3M���
3�,�<.��tkY;#�?��Ubo�(Ψ\j�PS��v$7����w��s�a�Sb�����r|N�Ae#���&7�<\�J�ͺқߨ6Bm��r`���t��1�5ҕ�~��A�q����y�<0&�N�	�_� 8e�d�]q���W��\��ð����Q�)5���: ����O�����R�s8*/qMYa0i��è���m�%X�<u�-?�eSȼ�P�M��!@���q��׮u�0�{6�8��~b~���^,*&�(���9�&� bNO�{��ޮ�vS
B�cy9��d���£�@�*"�8���3E���P���ȳ��D��*��g��*��3dK;��/���FZ��%4����Lgf]�׿�'���v�2+@A\(�U���z�{�^��<��:ɍ�����+Ր��3n@�
��%ƥ�L@��)��b�"����|ļ���}xk.>GV�}����2�JV)�����U��Wk�P�M���d؅bXj���>�x���٬A�D�a�4��zkx+����W�$1/�Q!�N��wb<�����X0��D������>S,���5'�J���x��+D���ϋP� 	�Uل��L��H.�{D�^@HT��4�x"Y��A��0WJO �&P�`Ꞇ�^s��N��G0��Z�V���p8 ��Cn���v ��K!�tx��Y�MG��vr�/�t3�}�O��3<�c�)<9+Ƒ���V9��ضz�1���˹���О�f@=a�T�#���~��/2_wu��+N��9��o1�&����v��od��	��/Oyu����I]
��Ӕ� WYJ��mVMZt��
���.�4�q��g���m�9���~�o�Q���ɐg��jL"tf���y9�:�ـ)q^)z?�������K1=��</�!=ʢ;x�G��8�6,$�O�����D�%��H/���x�������	!2�dƬ�c ��8]�,�����}HCH�0�B�$��L7KkP�R�9���"T���d�P���F�c�C��s��T�=
���[�����K#�n��jbE[ڸ����V_Z���@D���B>Nk�������A/ܧn2U�p�ͱًQ�������*��&i/)�*�~f	]e��+~~��s㭩ݠ���W Y���ýZ+�N�SV�����%A^d�Y)(��q��p��MD�5����3���u3�r����0�����/5�_*.�9�qy��Y���R�bo����\����=��T;-R�%��Q���f:�%�ْL��C����{�{�x����=����5�U��B=!�'ؼ�3�]�=7����w�5$I��c�ְ�T���߁��ң�S��V�tn��/DF��t$F�������(x��c
�Il�����D�r2�|��z��6W��c�_�He����'�m���7��Rr�)�^�? �2~G��_Px&]ȷ�E*2���P���f�.;�M,I��z��E�{`9{�fN9�^S�ȑ �߱E�M]y�8���$>d�Ӟ��t5�}��">�� ����{����Y��M�|�����.+�)���߁�"L\|G��ܓ�g�m�~�e_6c"�WR6�r���.B8���ۆ'n5��4�Q��
��d����g��A9�Ň�&��t�#�?'���H��s�~���D�B6V�"F-��"�y�|��3�)�V���+����d$0/���d>���M��_�^�F �`�F�m�#u�B'g����d��򋗾��<c�@u8C�X8��l
����p��&�b�����'��gR�4�V�0F�Ҭڠ�Xb����������V�B��;�@>���,��Hذi����eW}���u�Ox�hB��^/�F���M���$&�(MP���줓�>�:�hAo7��K�i���
g�����+�7�[b5��t����fᓒ�T��j*�P��	��3��1#{t�
�q���UgN3R�j���Ƣ��z?w�v��ι:�H�ʄ����W�p��@"*����3�b�w�Iݥ�����+w{K���Z���l2'vNG���ae{�گ/:U����J^����)���v��2��p��s��ڲ=�5w���t�c'3�v�5�ޮ~�JS�@�D�����\���T�/b4����%#�ⳮ �Ӧ�P�v��F��O�����w��E��h�:�!���򻕂�L�%�gu;��./���v[OO����+��pbN�����e	����� ��*����s�/^j5$͚�uK��Ww��r��2�D(�8/ �������L6'�����Kr.�|u_c�d��ܑ팠���dt,:湦tQ��&	v�����L�9OdJ�#)��/������
yJ�
a�I<�-�6��u��طUY9���2�T��eg�2g���(�����W�t+#�_����tŦ�0�9�`������5P�&�o5b -&����EG�#hl�+X��BFD��4�q�x^�m�O?�\�:O0�K�����Q��X5�T�$7�	�gP<o"F�G�����Ä3#g���������5b�YϹ��oտ��Qr�Q?����|��t%���`�ox���7h%'�O�q��ms4PÑY;��Gv��g�nm�>S��>�c�8+�9�b��>�K�r�"���ߥ�����_S�����S�������]r��m����I�ٽ��av�?w��65+E������T�8�ٛgeeO�Sv�l����%S�T=�P�{���IH�Y�����}w�N0lT�a�<#�F��<Jokb���k���鞲��١��]P�K&��m���!�3a�H�w�&
[,T^N&�Z�R�^���)���
<�j_G8��'�e	����2��5��=*������[��0��;�M��gd���w�OQ��]�R��������t)����\�
$�/.�З�S��+5�ɌH%�h��Ba���K�i�d� �Zਲ&�D���*y��>ʬt;�Ǵ�w��RV�	���9��s����[����D[(��#
ZW�����Q�claR̻_P��J��{�Uq�	{#]�F]�E�oҖ|[71�a-�rPbi�S�P��b�2��#�R]P��-�6歬22��c�V���� �y!PX�<��*��û�a�c�x��*�����Ӌ��u&�r�}���d�K�'���W-侁%d��`�M�=C�9����I/�G<�r��o�b�I��Z�뫻BRƂ6;�c�Ҿ�]���>Op�����7�ɻ ��m`��͋Y�Q7��|�F�,���J�9�w�+�l�u����/��Ѕ���1�~��-��R�L�r��fʆ�E$����=ԲV+�%����3��@��# M��M�^X�?��Ǘ��H@}O2�dΎ��{�GT��3E�+�M�'�u��mo����_a{��-
c��7�eNe@������\�Ɓ�ly�#���������/Ax%pݜL/�í&���12��2WC���Oږ��^C��AGK��_S��GT+n(��m(IR��)�'��.���l���t}�[�&sZ���`_7�Rn�6lL��*fV�B��m�t\w
j�c��y���Bc�4�����Эb0��s@3��8m~r�C�?=M��Ƀ��0YY�4D�P����9��<\y��1����j��.�i�^ڊ�Ճ��/�3��-\����o��հ"��"�լ,����eܢ_E��T�T�$�������Jϩ�7�g���ؤp�&�M����}�fI����YT���/�dGp��i����"
Y�@�7a@�	�R���B���u���y�n/���6�١�H-�`�y`?۞ƙ��m�y�T�~Ϝ����q�"Lt��gdS�����0��lIwʂli��AO������m[�F��eD�'\=���p�jS�>z�,�1���65�����fTӞ��F�v �fv�;����	,Ky8r�u�zUsW�������U(i|�BI�2d2d���bK�9�|D.�߯kQ�C��>���=#I�%���5(3��f}[��g�({$�1��oo�k^���]pq\��륌ƕJ | ϩk�<��s�@g���e;\��p�	��:/�&^�� Pϰ��}�I�Y��0�G�\��z'���"�����?k��tv:���Q��s���c��ӫ	�Xa6ueE�1��O���Я�Ϝ%tg�]m����zY[�>P4��=�%���w�i2�ybe�@$�C����DAlI�+I� �M���,��\b+�Sc,�(A����1'ќ-Hf	~g�����(Ӗ�U?N��B�������"����)�m?8s��&� ����ԐQ�V�PVGE�K�I�4��J�jvoKa�:����ۦL�7�[킧���_4�>�bg;d#론/+�	>8�j�R$�(�%�[�{�_8[b�d�[�9Ƹ{n���`3�h��v甋�����tf��*�����3�쏗�5o�IO�����j�"x��9m����.��+��M�y��6|E]	$�.�i1�)|-T�d���'��?����eɅlEo�~4�Ie��6ٝ�Ē>�(^R9��#��،��c��m>�$叄2}Lt͐�u��DxWNZu�&��)�Zꬓ��?+�^���%ݾ+���Q�o��C0�/=j�ގ"�a4�>}��ʑg������7بi3�,�س������Fe_�xF!�!��S��,Bؕ�ô�4�����+���H:I�q�N5?>�j��<9ʶ�?6�D��vB�.���S����o�?T΋��N����QJ�s�c	�]Ԫ@i�P����U: