XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��zH<{̿��ҳe����>{e��^ �᤬]��#XM�I�r�w}�Y�a輛|Ro�|\ͯ^��^��u��h�����r�
3_��&g~��j���7�wӄヸy�����o%�`T(�ķ��?ۥrx�&>�!H�/��F=�P�!���2e��6v�`�g��|�9���=�T_XVP=�2MW��Υ�mx�/\NztKG���Z�x���}�v�����J�ϸ�a������E��}�J�=�:?[�K����>]*)A\�{8�^�ä/�{ڦ��5%oP���{��09;��G���ZAR�D&%���V�WZhH.�Y�7��	9��^��If!�L�����D����wiz���A� ��a5P;W�V�6B�!����pq4`�;~7�u�*f���y�u1qi�0��I���S	3p?a�$�����]����sW5�i"9^޷��H�p�Y�vSctm���B�Z��h��[� �R�gք�?�H�!�a~jQ�Td��W�+�*>�l,!G��g%@��{bT��%��	v��m���-��Q�~/ہ4픹+�|�x����$��~�\�)���##�}i����+'��Щ��Q�B�ܝ�5�TZ�BF��O���Gx٪p���	����bG٥Ą���uu*j�ab&>|��TY��B�\vɂ)4�_8�*�;ʫ��Y~K����0K�X����r����|^<��-�`,A�H�&\bc�[,Lb2��x}D�q9��f��z1,�r�w�xݛpXlxVHYEB    3504     ca0�e)���ca��\TWˬ?%M/��z����#�\ �#�}Kg�5�0��i_�"T"�O�1��hM�� �M���AVԹ7�.ȵ="���ͽ��@�%}r�-����2��"�b�/ב��+eک�k��/k�K����d�K��ll+��Rc
��E���-��t=��}	N
�;�Q4��R��|��陡}��.u�1.�9����,��{!��1����M7�:KO���e����RҵzC��*���#��H9���d":K�4�caw�a4������n3XH�u<<_d衕�d���|�,�%U�O�JT35��N��3C� Tğ�kɿ;fH6X4��;�����:�����>�o[k�i�|��u1����]v�r��B�/L￯�A�x!Je<���L �,n�� N}�Aq�=}�^Ex��XA 6g�ITF�H����Qg���2��ˬRr�I炚���T˖���E���M(���^�.iD{Қ��[����y+ ���o��"�GN�-S�k8:|#��u�<���ڇ8�����Z����F���*�<�@ԉ�$��\h�NpI�c�%_ܑN��);$�E��8Z�tQ��I�.��>�u	���jt$�ݚ	�n��R��0Ö�C�:�pS�&f��m��Y`��{��r0��.�R�}����u�����S䲀]5'���Lv��YJm]�;��`p�� ��뮀"�:1$��q�{iO�j[�&�/�~jϐ���.���Ec������g	%���X5ZV��x�����|�6F���9f�ލ�r�8j����΄IXrԱ|��Y�qu=ղZB�A�۸�Ţ�,�~쉋�ӌ\V؏B�~�V۝^z��E��y��v)E��JY|o�T�:-wg���Jھ����]�n�ܜ��^A��J8D�1>�^ڤ	C�
����t4���`}3�p����e�7��OcZ)�qp!�Q�?�r,� Pq�����BǕ�X�%�5g�~�}�Q2u���2�V�o?A�ӱ��1<#-� ���)�io���=l��d�7q2��1Q����Ԗ.,|ŉ�/o�LJ7�I�Ha{9��Ck����Q��@}��jJ���$�R#R>�>���)�KQa�4^���{��Q%W����1���aC�O��p�[l�ds�AK���ku�yڙ��[@���d�*��k�,cel�bCY!/ma��\.o�%"��~ ]ew�ӡ��G����P������?�(�$����Ge�w��'��\m�Q�`��-���u�|
�=?k{���@����D��fUJ�]�8�qc����7�g>b����Z]����ȁ���{��P�:C��uu���W�2�;�)-D�S�of� �b�E�Q��ܢ�)����Xn��,����R|�+凢�$eS�8�<��>�eyA^��xP�Q��������n������#�>�*���	��W�J#i�&�̧���Q�ëT��p�;�%_d����,�a1^���Y6}�(}d'��X�$������;(63������WBg7�
�=C�Ѥ�.k���a�{�7�o���%J���,M���F5߮I
|y�o��Gs�m��6�I��_��e=2�e��q!;��܂�L�Q���������ز�%-������e˔��К�G=Y��N;à�Jq��ڤg�8�Ё�ؕa�m%4����GI\�#/��}�]���g��@깩�&��ۗ�3��ϗ���0�2D7�4A:��"�)F�mF����
�����#M"����_��~�y5L���$��Z�E��j@�XQԫIw@x�#~��8�<�;k�+ �'�#��2�y�݀��E/���k��t�N樋�&8K�VC���d�oQ��0B�R�N-�[(|���SS桐�������3��*�ӂ�ayL����z�K�1����?Z֟������)���G���gc�5��/�#�U���ͥ�k��c��Yz�~O� #�X���^�U� YS���_��:���lܸ~+����G��`��G�~��Р����f��_m�ڑh1�����#]���|^�CQ�)`�n�ǅ�;$�S��%�W�#�A:T��g��Gr�m��$8�k��A���|a���N0��?��nta�	d`!P�R����#���%���\�:fLJ\�����d)l5�,Y�cDMDj�
� )�~��q�P�ǘ6muz�90<4_��䶢����IqX��g�Ӵ�������u���ț�.����"x�5�0X?��׶���f'$�3"�c~�}Ð���D�����DA4Z�?��
�8C�_�}0��;*��%�A�!%#ӊ[�u���\
_)���Y�>�'��Th۱I�
�R
�d�������n�FJG.,��ixN�m���ᛊ躞�D�-3��m�Rz�
��[/l
�m��YF7�5�ȶw9<���O��>���&���D��g'�5d[s��I1����`��1x,x]�A��Z���1!(ȑ��W �զ���p�}�O�첐�ɎEJ/=�n�
��nr��c�/�Rzu��k�c�A�&�f䗀$�	�R	�J�,����LA�4P?�6c0n�ź�_����ҭ�Qʠ�Hשc��>�NCݳ�Uw��q�QYJ�QjC6�:a�h�'χ�q{Ψm)�S�ߧ�D1v��>��?+�����'?���2��d(��4��
M����U��4��xZG������[��H��ڡK҄~2�
]����_bw�HV�l����y��We�D�|}@q朲�[F����8
/G�Z9�[�#�"D
�����S%A&���Y��M.���=�e.��@�֙���L��{�^Dkj��T���5U��8��]l�!t�����[|��c�Ñ�g�A�f|p���+�k�Jj���bH���ײ5�/
Fd�.������mf`� B��)�P�k#2�/-q��Aq��%d��޼hya"(?�G����7[j=B]��֢�~���ׇ�C����S��7���[� ��N���R����ϗs9�	L<9w�twC�ck-��/\,k�z����8;Z�>�� rf�|�9>�[�$�ҕq�.AF��b�r�5�7�o�-CN}<v��X�B7�\�~ܤ~��Q�$l�#!�<#s�iS�f*d���A��$�;{��6P{�c�u`