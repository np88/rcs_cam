XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����"���<�L�9�v����X��W��1h���,_��X�_|G�����2&��' :mU�Cfh4v��\�\�m��zdߑ��"���nY�}�Si�.^8�L�>jTa`�.h�Ҳ!4�>����J���C��Q�^���/|�a�id���y�RF��A��������׵2W��|F銺V�R/�*-,U�N�8��j5�L�gqx?�� v��+����v�,�QStzrR��8>5�]�*�N������,��%��� �
�������oy�g�������+u�ſ��
��G�m�\=��rN�)��k���#X�F�� �,����D�uC�S������8�P��0K��@��X�T�M&�Pu����3c:��vG1�X&��3f�pJ��̘Sq��E~��:�X
�t�ϣ/![��Y�:��i��&kAi�C���A����{n��K$i���D츿x&H^��3�/�����ϻ�$ܐ19�y�|ʑ�u[�X�����-��J
�ǲ8/�_����73��:�#/�d|j��D��� ��/�Q�b5e���'<l�����D+x�ԩ��1_fw��患ᤗ���G��$�.,*ESJ��^���M��I�!R�f�u�����(�J��M�k@G�QC�WQ��ϥ��A���r,�8yPN�e!׍N1�שŠ��=r0r�뉬2�y������i�²�9�9�>C�Í���t*� G<L~Wna�#�x6�Yʝ�X>�+n�g�u�%ZRXlxVHYEB    4fdd    1090�.��Kx-�t��j�P�i4�/s�=%��C�������3y�߮U�G�*��H ���@v`��L���/�	"|�\�e��L�P\���|ssLp�s^�D�[~N���-���ڻΖu 
U��k��T�
�Zm���\��+ah��'�΀�����B����i~�W��z��u?&t��w~��'�; %�N����SR�X���4����Yn�G#f�+,xx�
�Kn�M�E>�s��M��b�r��и�_�1����������lC-dF}S6����~c������D M��;��P^[@���i{�xToO'0P߄��ζ߂��~O���!�YI]��WNn{�� R��A�X�L��ނLDVm��#�(iP:f?
�&�.	�2�<��	ځ8d��2�����v�	u���WWX/W�	':�
6|��wp�ğ$ {�nȐ�'h!�T3�3w��,�Z���(��A��w��-X�7��>��y퓽_ <l ��z�Bv�r�X���5|�E�l�Lc��H���a�{w�b����ҩxq�\a��=��})��l�2�M����u��j6�5�c �4���H�O���*������
�b|EW6�A��X�T�>����KCZb�'��OG�N�eu�	��vQSi�?wW���2�I������!顓�Hg�i���n�����b�c�`�V�l�������JxQZ�\�����\��c�������C�eaM�m�wgC@��F�e���934��N�5�7�� ���0yL�;z ~�d�"��3�}����Z�0l`$_���Vό�����=����;�N#���Dp�$3�M�9�A�[��+O�BR&h����;���u��4tN$��{K��Ǥ��ydO��K�@nU3��Usfv��f���y���蕟D��T�s�?�>�i���܎������x���@�w/�@���\6ϰ��ަO*Q8�Zn/�]�$��Z��/˪� yً����x�����P! �ays�Ul�(س٥4�ڃ�vV��H�#N\_J0�-�A#������=����J���K�[�Ē?����~��㸷A����h/����
At�]<'��9
-&�ҾQ.�� �U��OP���=�;۳��p2\�ْ��?�'�z�D�
�����)���8�Z�{Tȉ���A�̠̮�������xd%��<"�?��>�-'�Al˻�ԕǂ��n �W�t�_��$�;h`L
��n��0�;$�����1���ļ�-j�֥�P���k�2�t�0r;F{h�ԙ��}�������?{z���K�A�ɽ�_
=x���&'S���Qz@$+�
l���|�
<4��[A529�qo��4u�g4'����\���HBYL���g>��U,��z���M�/�0�1�Ukr+Tܷ�����0��BO+1ˡd �{��k�H�HdH[� �tb)���������c����Bb����2�r��;�k϶^<�:1QG��P�"��_$%�T��/<V>տ����F1�)���3n	Q���u�1̶7�2�c�$����0�b�B]3M���K;��{���b�#X�Sx�b�Y2���Q �¿��ȃŭ!��1�&ߚ�vxy���Q�u#ܒѪ��q���ڲE���l��*�x��B
#�d�ޙ:���:X�h�������C�S�WJOVLBh�Q7�!{��9A�M�^J�� �<�h]bg(�
�/�j�e�Z����	B$R`Ϧ���a֬f+�'M����ԁ�`�O��B��]�e���g�M�#x);�	��d��cs�=�dM�ot�	]�g��Z �:��G�]�*��WUP��*��)�D?e�bZ�`���n�j�5Өq��/݂�HS��[ac�)�VxjT6���\y�Mֿ7�$�\+(�?{�ȾSx�����b\������]T{u(�������=
�ؗ����h�T����{�u���dɰ�r���U�>�j;f3|�1�T�kr��/כV��<�V���2O����t�^�^����
x*r�J3Ĉ��%�-h��{�俙t�5UP����((h���ꖚN�)��`���4"�O�!����N��۳��۷�/v"T-�s�Gq��a���/���u5:���[1}�i�N����:bARX`=^�d�8P�^:@]\��V�p��~��$�3=�پtZ'E��F�'���es�Z�29�r�s�]�>A�c�^׼k�.HnT�1p_�AYTo�y�����t�z�$(�}��T�^�YХap�D�wAbLVQ<�iZ����p̶i#�W9�%u�^���.����Ns�1��ARG+O?��a��`i:^��
F��>3��/�EX��9���g��"W )'�H�Qdl��E�t���!�
�Nr�g،�B�`	�m�7�Z�D�ޫY�J����m�!D&b�v���r)�� �g�v|4�
3"��-i�o"�c��%��k|��>&!~�p��� _*��n�?������&6������{*���.G� I���qr�܆� }�. ��V�cC�n���s��n��
�ɝK��0�\�U5|Q@����3C_���`��ҟY����'q��0�L�U[���Q�O���=*����-;���
{%~~,��n��ԫ+M��\���OԹ�C��w�[��~6UʹQh2��[��F���Pk�}�"�j{�0�^2s���M/~j��ʆ�����jA��'��Of�2�{b���QAż�X9h��1
�?��*R�]7�N�����Ƞ�\pU��(#e���+a�R���Q8�c%+�<^䯻�;%'�Mz�|�1�7����@�ѭ��xE"����(��Ea'Hb� V�rO\ ۃ�*��u�8��x�|q᭍�&�fcO0���9?`�}�c�`�c2�Z`�I���a+��k4�3v�������wHC.�5�V��1��WP��~�q�='+����	-�Y<�b�s
7|����)�8���E}1fbf&��E2paG�ÅO���KJ}�
r�	��4 ��f	3?%B�w }���8Ħ:�d���^��rˋ��H�V%�\�G-��!����(H�+_������|�w5(ۿS���<
�#/���ݣ��}Q?[�g�wS��V��@B��ݨ�NV��I��'��H_EE8cfԩ��c�^� ���x��p�u�m1�X�d?�J �BRb�l!�`u*����A��-k�5�y	4Q�}?ꓺ!iy���f:�K!%�V���zŁ��Y�
�֧��.�%����?�p��g�F2LzF��xڌ*$�v�.�G.�gZ	�����z$6��\����{Pe!T�$t'c���L��y�]�E+x/�Bbo>��*�|��;%�;q��7�A��j�Ȣx�g�T���UvJ{��笇��pI��
+�M�p� ��.R���8x]`��U�2��d!��j�=��c�Qr_�+���4cp(n�W�$]������twC��0��vP{��j��ra���Ŋ��&-� �ڥ�����2�TT ���C�;ȃ�u'
�#���C��_��hs�$�J�m�m�^~2��=��@�(����f/���V3o����J��'�O��Ò��|1�/8�4��#����;}���{���	5��W:�(Rc�$B�S9��?r���H�d��h2���I�P�U~aw��i(�2�9���W'i����ӢB�S���0~Y�̳�>$��`�yVYTh����`qԋ|�:����D3���c:+��얋*�}N�����]LY#9EPn$W��˘�,�p��ɿ��%���M����Gu�R�8/KN<�U�V�n'+}*�7ާ��a9�)�:��H:�%�2�68ҩ4������me��At#���~W>l�~�W�Em�l�g�� HUnT>�T�
�к��������>���-H3��W�s�����k��_k)��1��s��	h�%e�O�+��U$m�hO�����L�`�`�0�o�A-�Q��!fE>É�6��'������d<9�4ߙ�r�m��~��B(��W�ϤzDa��8��Rt���#��T�a�i��\L