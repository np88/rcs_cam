XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����dQ��
��`�r��3?���o�E0��攦��H95�ݱ�,`�bt�4B�Y&<�����R%0�!@�~�B��z���3��k��R���2��	�鲸kdԈ���kHlL����������T
J=���)0~^��O�����Q�$�F:"Lɡ
����;���k�-�ve��ђA:�V� �ܫ"��[��(��`|��SI�L�������EoPi� �3����/v)��8�6�_����$A�ό�c����_7���;H�Ò�,�᪒���f��۠������$�D!���ܿ��W��rf�Y�ܐD3v+��4!�$ѱ�������-S�B�Njg_�B��{�^�*q��I�Pq���/+��B��<��p��)>PZ�K ��A`��6~�T}�Y����UmN[hq�ϋ�6��C��(���+2�GS�k�3u�KA&��>����`�a~m����!�)��H;�L���������{1��	�\��X�Z�Bd��Uch��B�jp�K����*��u��l[+e�'����E��d4�B&-��j�~�5Y��R����d�5u<-(j ��'�ս��Z�/U�W�H�S�15�8U\���嵦?І��芘cb�曚��'t&Ҿe��������4F� βy`����bת ����l��v���a5��k/�no����:���]c�����m� _��Ruv��������>��E?��Zn���qy��8,<�XlxVHYEB    4a8c     ee0{^0����e_�b{	R���n26o+_��1U��yT��FW&�V��7��-�>
�z,1c�G㻝KV�s�}ѹgd�Ӯ\���k|x��9��Ά)��=�M�� q�>ͮ���G���`�;�H.ܦ�W_PƵ��Z�<{����(囐)Ԛeڭ{b��#6e�*�Ni�e!n?�1��x ��SƾD���PjP��p�ẍug�v�F!�A��6h�dyEإ���90e넇��m��ws-�r��o�V�tć��K ��o��XX��o������gc���[���z��V!���DĘ0m�C
^��ã�.�X״9�#��N��q'�@�U�5f"��bu��j��.{�|#�mf�oL'�~�na��� �����m�f4�F�g]���)PTQ呿RJs4Z0Q��`���W�+!�F>3��㐿YM�����Q���6:+J��;��1q�Y����`C�H�ګ�Ҵ��,!#�����/ø�B#H? ,����Z.:�+�L�Xp�3L��M e�ZK&�&6����nF@}��,q$�/�LY�~��a���"�k1��{嘳a���:�ؾAn/{Y2/�ңԐt�pf�LR�\y1��N��Ӻ �F\�d��w怘�������3��q��y?�.{aC��Sf�u��׉���D����0�N�,4���T���d�� ��/����틎 "n*@ߏ�1B�;{_���'�q|%e��Ûm&֡ݓ��~w���|=�$��o�}Ď�j���d���(�Jyo\}ӵWh��%�g���.%����Ga��t�8���85��ђƃA���n���F�χb@�4D��y����U��7���f\�Ẕ��;BO"�t��dg欵�� پ�ɾ���A	�Y��g�b? c�����?����ҿ"J"��nC��_ee+�ѕ��K~�fv�J�-��qkM�HG�jy��1S����f�'�
�rNzs�i*$�'<PB�{#6$�t��*�r]W
m3n"ͥcG#�Y1��bB�42�7�����?���c&X�c�%���*�D�o�O��	���J�I��_���È�8��ձ_ZQ���1���X�f�df��t�k�^~�)y�%̼�G�����Y3F�֦��xD���d���7?�����:�88�3)Z�.�Ɣ`1��0*�K��������T��	�j�}��3�f�
f�J�%w�Y\��*��Xz^s�W�U���į�Jx�;u�c2�h��:~�h�<i�D5y�UE��?�T6:�f�צ5;��pݛI��g;,B������*83|�4�-mi�{W6��1��͔ dz������_GC�?O�S�mK	����y�#\�9a�
���t��%��U���Gg�xDMNbc�oe��r���dA���Sʇ���z��*<G"k�����c�3�j:�EGH�s��MoB9���,�S��,0�e��b�0�Λ��:S�Zc��$�>�H��q��xn���+������ǚ�Lh�!$qk�^>��!m��`����֟�
�>���q	alH��"3�E����U��I
2@Y>n��T��o�0�aE־��K��*ro��t݊��Ι�y\�k��lf-o��;�e� \V��am��(��t��Ȋ��>��ה�����׭ֻC��"� �+�(����ܭ/��FaP jd}g�!5֪�GdӞ<u.u����u�GI�|B������e��2oH@(vB�͏N�ޭ� �q�(1&l��ǀ"P�&�]�K�#LȘ�k$(0��X7���Ѹ��P�i�/zHr7�!�����p=��߾����j�����ws����4T79�'�tyo�t3ڸ�������7�:J3�oA/x����@�%걞�I0������^2jYf��F�z+b���S�1>��M]#���>6x\����oX��B�������O�VL��<���<�5Ο� ����+tGeY�yx=�y�0��-1���(�i����d���x�5j����5�:��~�#l���^��oPtLR]I�C��?��@L�p��>�(��:�%��}���or�E2�6D����ᤨ%T&T��h�:B�R}$�K�c�ݏZ%��^D��������+���R�����cU]���9�\H~!�/������K����7���O�<1~���rp��E���6�"F���^ ߶�.J댫��\%�tK2�+$扗|��E,`��3��D�X�p��4Jp@���fhMe�{NO������^ ������>�ezq�HR�B�SO�o��X��AY,E���W�u^��y��@K?�ia�.�f��)A+܊J�*�&B�G�O*���D��5@�[�&>a[Rю}v*m:�ck�祼���>�־�67���7�����J]V�a�}�C5_/Ҹ�.I��Z]��?��V�	n���9#���4\$�2V�u�0ˤ�����ô�8�Je%ݍ�8����4�ͼ(lNw�71�ʊ	^��T�R�`0J�V�N��䏡s�U�L��.1l�a�G�)��[�)��7ԍ69	����cV�7���p�*�Sϐ���<N��i�W���X<NN#@�/!kaz;7��~��o�Þ��E�R����G�WS�递��T6�Sr��8�0��������ߋƃ)�M�������`K��������P�HR33'!)���!�|�+a-�S����Ƹ*��jfդ:FjXk�
����3���5����묖�)�*�=��H�"�()/��]S!j$�X��2����I�m�BT��pI09�F�e�݀S��8�8^��,�vA�q\S�.���C��5 9o�oG]-iGZ����?�����\���)���(>�G���3 A��q�i�m�B�׺�{#�~$�ޥ8�s���I���C5��j��1�G�&��Z�y�D2Q{��;f�
aA��d�@fC��[�a��X�ZM�j���ɗ��\2�Z�E�~L���qo�:_X[6��s!�w�*R�7���՚�f��VX�!H�m����С��Z�̤Y�4 FaӲ�޹�o�m�(��"ɿZ����Ӯ����эc'�oizs�e�0�i|y�Q�L�[m��޿������`C�w�E�ɻF��%����QF�젵t쓉�El���L�Æ�_s``SG ��*�"�{�DX>  0�9Ad�d�J����@��s�MĶ���j�\3/v�2E��KZ
j��ٕ8��i�{e_���#�.�7H6��^3_.jp��r�s�EjN��:�D���"�
��(��T%T���\� � n3@��� �$���L�W��'5���\:���Y�uB&�q�����RA�-F��( �U����i�UÞ+����s#�4[ǖ�����`�#͎���e(%����E�8�N�y3��죥�(�����U��A7�6qIV� Wr&¥]��-+DG���Q�i/J��G��qx�����z~��@	p�jϑdU��K� ��ҋn�<3���jE���0��z��*��'�7�,r��n(�!t1I�E��Y����%]d��Q�i��Q�F����E�P�[^�*M��8�@ñ��z��uò�zw��x��3�wg����~���+Y��"�:%N�2Nb�kG&��#tŠ߆'[uy��2N�GXY��4,�&D��$��	�7Я�s����y�b�*��\�t���9�҅�6�K0n�,C�