XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��b�v8�'���Y��5�]e�Dk� ��ؚ{ava̓�̬�(�y&a�i̡�[�9�6��n�*��&�Lata#ǓȋM+߷$}.�eM>���:���ʕ*�~oG��ǲ�&��S���9�2��q�a��D䥶������l}1ˡ`�P;P�?F�|8�lL�5���dK��,T��h��(��53�eG�re���hn���7%̱?赢���4�>+�Z���
�M�є����Ij�r9Cwᤛ�"T��aMl��w����@J��K!%�D���U������%b���h�u���螇�F6J���Ȋɂ����vf�ec>�)�L�(e��k�#�~�m���n/��\��t߅��
�j0���tz�bڌrXB{�n��)�7�lu���A�S�7yܜ������_��B�#�1Z�8�v�/}�����m�L!����hX�cj�F������Jf*r�+rZV�G�Q�-�(�
����ߟ���j���'�ثhb~�=A��o� R��+&
��Y�$��0�j�9\�yc����i�q	��d�X���ma���hs*9Q���`~�|�����A�6��6'<�9�� ���F>hw�r#����s��}OQ�j��U$ؑ�nz�O�h��r�`���D#���$Ї����p7�G��V�b1�:l�F���e�Z	'�>(J*T'N����{/���F���C,,@��\��N�`�O� k�����Gڊ���{G�s��1�TW8#�х�?/i)�7XlxVHYEB    1ce4     9e0ee�]��4�=�`��h"�{�Ӷ�p(f>=%��9d6�e���tU$-�.��pty���h�M3a[�����pQ^��n�c�s��̝s�?�������~����e����|��J˚�XZ�(�z��Io�w��!�Vqu�y;�TXMʶc� �;�qSΥi�E���-��NK��c�$�� (��M�n2k�o�2�5�|.sq⑵�}22�[ھ�]�`<�jK�ݹ�'sk����%�\�J��oG���AY��'�G���o�m�G���s��c�3�Msѓ�5j�4j�������~�잦S-���K!�L�_d[oYo,�=	�hO���N���0�m�������o%�4t�$~Zc3��S��{g��kl�?Y�r���Il������T���|�D����ѱ�E����a�O��kN�� ��K\a���\�r�\�w�T���P�5Xj&q�]Y�*�z���F�,(����a�lä�=�o�
�fN{,�i"o�8,������r� W��0�{w��Ғ�Q����v&�/Z�h'�=�����k�ςE�_(}����*Xbz?k�*��;������>��;��m4p��iB7�d"ue�ԓ���Y�5�*lyᨭ�lX�c,^+7%/���VA��.��HY��ꈂͽ��W�3��Q���ƃ��oL�a�ۊ�WWd�����sd2��ʧis�!�K<(�?a-~GI�y�Z�[»y�3�,�;������{K�����7�t�zW���]����sQ�ຍ��K�ɨ�8�>SN`��gs/*�S�l.y ��-˾S6p�겞�~�e�u��~=�1ʀoM�O A�0��K��uHI���c�%]@L�)�׹�f���K�o�$��uS>;Pd��M��}�`j�I�U\&�c��"��`K�CF\�ߩ�&e���K���D�v����C��~fYk��^@l%M�N�%�j���Ŋ��8���IbȒ'*�5ty	޺Dv11�N3ϗ�.І��過)��\�s�n�DZ>�dKU :!Kˡ���D?����BG�~O���q����0.5��#s��K$�#6�M��[3$�� ;:�F��}R��]�!�`���b?��P�,$ԅ=�3��;C=�{�A�4���2sm��]��+�;z:�N���N#��E��=�y�pLJ�V���D;æ{�U]m�毤�@Oۂ���(%���E<�q3@���=��e(>JP;�c�_G�K_��Xy����`�-���nb��}�u��Ws�����W �^���:��{oglc�x���9��t�B閷Gt��)�Y1�̷N�����`\f��!a����������}�����@�+����,|�d��58isIdV��\�����M	|-��%����vgA�$����z�����P�:yOj��U�9o��$����V'�����S�l!5|�gGX�2�Q{����_V�$�|h]��msU�6���s�x�4�s�3x��{��=Lup�g�U�=�n���@<���e��n����S��h&W�L$p��br�|��ޓ����;�yx��/�)r��2��a��Fk�l�2N�2P�S��T���ҝ�v�\Ɗ.pyp�\���ZN86�/�l�n{*������`'�8���m��g�mx�,��]AtB��^��[���*\�����*�5Pr[
�`�X�F�k��>r�J��
"@�vOظ]13��Ήw���5���~�(F��a[["pM�(�&��,����6���80�Sc�s��K���W�U��*�D<+S>��i�{[�}��rq��O�,ۖ����LRp����)ߐ&���YQ~�h$A�itd��ez&��A
޲�b�&tČ֝������I�W�X ��D:W���Z����7�B�`F��\9eN�|MS1��۰m*�PJb3RL��9"	�\-��-�$��l��R������Ji�@e/ρ|�#qHHf�R��d��}=��T�D�Cv!�u��Q�1$4F.�\�Θ�TLo(,C�3������{}���7���{�����{ˢ����2�Q���1p]��!m�PB���cV�[b��%d��|9)U�g���̭ì�K�Q��6�0-� �˂�SU7m��|�/��f{�˂�i.$.�B��"�:�i5�D�_�k��4��e�� �Q�o�YL�>�����ÿ]���b�S��5o�����h�4�-�����=~�e���.ҩ�;�Hb��_��&�	�T(�Ɔ0]�q���%K59a�2̩���L�`_���:��� ����¸�������"�����u+<f�w�U�g�����+��0l;�,��⡂E���ƫ7W$�P�4Om�3�J�਋��>0'���d��F�-�)�VQ ����Li�������8�_�|)g��� �\�E�a�>�c�x���tӉʟ�����y�q���W4G���w��'#�2j
l