XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��6�wf:g�0�u���Ni�C��Z|90>�D�>�H-�s8'l|�Ia$Ķ~�B�v&�F(�R��bD��|�ut��HE�H���R�D,�U	&�y�MDک�)W�pa��� Z��*�%���j��s0�"�����F&�.n	k��l���:�|#(���xx�V�~�%�Jnnk�_(a�WXYLqd�g���*"��W�q��i
�I�-�q�H�|C���f�b�_S��jx��C��b��d�b"×�1�5���ޣDuH\+d��e�@��wx��"��~g�0�/��06��mB�ײ���+Cb����O����g�\O%�,Q�8]-y�/gjJb7q����R���\r�^�^�y��"�-��\�}����?����y*�1�d�7������lO�x`��%���қ,�(>/}*�}����� \T;|)B��L3���������L��t���v=�����?���7��c@J�ma�w��{���Iv ����%����������Ŗ��B�Yk�r����Z�~0W�v��#300a�Wn�K<Ogz��XC�j��9���������./��1��P/�A�@���Ə3�c%�U%��[�uF��Ψ���C���1�ޟ��qi��Loku�)�d�bk��Z��VĦG-͞���1"Xj�\ܚ`��/̌���j[{LѺ%����h��@�� 7�sj�B��s%����)��t��#\&w���P�����fڸ�l��H#��km�y�WFX���rU�5T��ے̈XlxVHYEB    1427     840dw���P0���)8d%��?��H[2�vL��Xu������ES�����%��&3.!�)�e�5qb��]/���ƼI�mU��U���0>y?1��X
nDj�����-Jq�r�����a�3��0'+ 3iŋ���*����Y���Q�L�5�����5NeR-G�� �[�Fb��3�2���G��_*`)Â�ɺɡ)1q0,��ܕW��ߜk�lNc��<X5}1�\�qU��) �f����:*@߿ ��J���|r(��B�����*��:�d�B}��1S��q�Q*�|��*�j�9�YX��?C3��s�J���.�Uu-ϑR�L\֋e�Mʃ��u��g�rߙZ�b�q	_�A���B��/ա׼���8�� -���'֜�B��H���<=6�z'HؠZ$x:pU��Yv��@�ʬ���Ze���y�j,�9��c�v�!�"m֢�Utr�Ofa�sE��w���֑#��US��}=F��*��۹�\��w?~����Qߑ�� }��=��6�T����_�4h����k����
ͬ��ڍ��Cb�����T�
�$�<�X�7P;��]=��L�'9Jr�#���tr�vON���0g���/��U��v ���:�6`8w���!�vG֭;Q]^�`n�ނ)��9�.	�bM�H73s�^U#��G�(
�?�Bϯ�����j�X�,]ڄX�}�U��6+��S�o��g8��s�,�z�c%!	1VY���y��0C�����.�2A��e  e�z�;�-�.��$cr6��Y/�6� v��"t��!���/���gl�
��L�t�ԧ���.}�-����w����n� ��+D���~����9���b�ӷ�Qw�5H=��kj%�C?{p�Q8��u;} �s����U��x���I��������%�D5c�p�Ѵ�5�O��O�]�@����m��v�bh� 0_����˨-���FXn�s��|S���)]�#��8������>�V-�t�P%�'_�+�L#�(\��n0��� �c���P�:ۑ���:�o�܁�19�� ~zA ��ͷu^Z���TП�)�(ҫLVZ�>K�L��+��ͅ兵����u��~����W4���z�m�qN�CEw�0|Loy�����>���7粟�"B��
5��$���=�h|�0�.k7i/H������7��K���SFX-�é�֩'���E�
�iұIN`X��^B���$UW�C���J~�?�X��y'G{��o��n� �[�-�)O�\�ɽ⽏O��� �K(Ƅ�G��!�Q�^�F8��$��k[Tu���!���m���
�J�p�<����'~y�dh�J��Q�M�%���4���,ͮ���/OCW��N��>������ɕXtSܙ/��"&��B��)���$@xz��x����p��J��]y�Нb/�]ԝy����6�c� [�z�=2�t������2~2.�].�'	I!E�r֑�����FJ�Y��eߙk��9��U����fڰ؍�����AY^���W*�o覐j�oH�$����]Oov�w��O;�*kd�"���Q�Y��&�����L�8���p��Y�59{��QJ�V`��ON��3n�v�t��k.o�����(3l��qR���CM;�1�t�`m��D%L��P*d���>k>�t0��6�"�g���kO�e�%CE�[�}�{�ߵ��	���z|K�L�D$�y��[Z��D�'����r�O���a{��'_�8n'��>��*~�ݡ�(X�X��m4�\{��Wj���,@�6y�3�+[,��e��iz��]?�6�G(�Dq��+�l<��+�ե�k]8���]�| ��%������k��PO�q�N`�#��Ӥ�>wP��K;����2�[�@��Հ7�:z�(���j�f�����͆D����gv��/�k;4J-��V$�sK�P�>��á1�ə�m.�������#O�7�����wd��+����+���w��S��{��M��`!8�(�+�0�'p4!�}d��=i��4��!�fGvn