XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ťc�E���N�*	�,Υ��J.�|�Yst� \j��/8ffA�\�F_R$0c�~6ƻ�:��q�i:o�r�_J�h�5�z�~���a<��࣭�v�~��xq�[p��3ȟ��b�饶黦��sk��'�;fQ��Ϣ�|�P��^a��n�߃K�|��dJ�ʄ�)U��ۆr�v^<^���2a�lA)jKF�4�
d^��⼼�ss��i�l,)Ԇ�Rѯ��NҾ��o_,r�ʜ�n9�E
5#�gXX��^0̘�R":����U��gա���^�?D��jXl�ǲ��h8�������ѵ�{f��&����.���r����ȓ��0����o�[�W�i
��ji����Ql��4�(��&��5~����D5���,L���!lq�΂�/�G��o�D�E��p��#���д�,�o�A���L���K�H��[�K��RK�tJ[��CZ�P��iX��4�_q�T}����$�v� ����_���`�bR�V@�1LM�W:�����Z_y����)����~����l�Ȱ��N>!-���X�|��!S�}��!�w��n�/)�ҁ�빵�ź�٤Ǳ� dy��dH^�;\s!2E�������湺�7x9�%穻��1Ci����7�5<�s�<%~�x2���S)�C��T}ꂾ�o����"��,���|��X��S�*8���}vPj{8��;�Aft��+�>՝+�.�f}�'�9M�E�-�#XlxVHYEB    fa00    1ca0���X��1���H���"�n�� ��zf�Bv�{ij��-_��@�c����H';�����4O��%�/�W�%2��)d!�WKnѣ��&+�#���丏(������l��M��U��۫,8��"$f+��WB����G���ץlr��IA�Qu�
�ϯ	�lH�Ծ!��z�l5��?,�e��E�)����E�ꌖ2@��`wl6��a�̃���Ӣ�J���.,~��T�ah&v}8�~��&�s}$B�`�a��\����=�4���W��:���@ X"IM�l�H=�P��)7*
�A��+�����a���q��r�� �d�_�vXm�q���%7��z���6r�7��z�2�nsB��R��P��9���/7�d&lu���7qnCd���.0L������ԗ�A�Ûj�H��n�%rj}��Xݣ]�_,$ϲ�������7�;��k��9��<�Hш�ԯ���а�����(s�ӿ|9_4<���"J�z�<K�C�>���!�c��r�vK-�ڙO�y��!�$��p��;?ڀm R���ơcJ%���C�G��w��Q��	�a�ʃ#le!�~z���1oC�I�:��t�ȳ��@�h7ˀ}�����r�qX;$~�L,4\��u���HȒ6���,L��<v1vt�ǰL)ޣ��1���;5n�Q�վ�_��(��yI����W[�R��Fw�|��<���X͇sC�c�Y�ma�yhH��s:����<�XKh�����8d�%;"c4�% ���U�H�V�%:ԂlC���Ž΅Q�w6��'k��ߟ�̱���˓�)t������w6��e�D�I����v��%��{�`������$��)݌S�ҕh�n�1�߻[꧉���é�����hKH*�K앯(r*-��6��;kԔFi��
���j3fC���Ҿ6���+��_�<M�t����c>j(�o���_��^)%�*�9�9ܥX0赓�
*Q0ĭ�x25pS���fOCԳ�B��C;�lM��^.9�K�#�}浇�?V�GÈ�:U����-�JN+������/��or�~�������7,\��5��B&��$sdS�@�5�'_Ps��, y�c�hDn�Rs���%"Z∀�
a#'6�h���~YS�!5�\$U��v�/ x����X�0�T��'x�ko��9s\>4��.��j���ۮ��.Eog��O+��i���T��A���L���$'�@� �����@��}}>jRF���,hF�1|�Y|D��Xa�����{r6��Ö������Pk �b�aW��a�f�n�L�G��V? h�w)��گ6f^��c;K�@Ρ��
�wC����D�P�.6�'�F�:0� �,���F�,]�XA��9 �oP�>����=��+MX~>c�I���B�9(N��6��ۤ��gkp�<|Of]j��ʩ�
N6:c�DI�%��2���KB�/j�l+=i�<��Ǜ��c�2�|����N	6�y��n_I)��g��(KNȳ�<��zj$�
L]�E�7����g�vJ��f����~C����g�u?��(q�Yq����+�#PD�W���%@ƻ�*�����*"b�HX-�W� v�U`&X7�X]Jܷ>ˉG�N:,'��p�y������t�̿n.ؾtG5��E�����-�L֥��Y���6d&���؍zg�K��Cn0��ֻ�0�.�%�X�X�s	 ��Azn�]q�s5�8�zXy)�,�n�/v�`�����>Ͳ��Փ�kHQɣ�`l�y�"�\EC�a4<\���="�yj�A&�n��m��J\Y���~ ��+���N�q�n����u۷F�Vu�[�Mؗ�%]c��Q3{8u�л�Wᐏ�N'�'R>T�\��<��9u������q@D��΅kY�l�+%��*�V�����r2����ݷsX���>;�����c^�6O��C�ݍ�*ҕ��͈M��@������L�D���� ��&��)���!EuJQ��j�D��=Sh}��5�f�O�.x8ǖ�/a�u�rvoT'&��1a3%1	�p���C2I��wl�H�qi���eT��_/�r�ˣ���HG3*�XL��m��k��7�_���ꉥ�{V���=z�;&R�x�]��=$i���[�e��;�O�_!RB^��םZ�I]��X�<����DO��`j�Q��n�faQ���������M(멭��_i�A#�å��t���D�gKt���l���s�͒D�Jy_���������W&�i;*Eh�m��V�S����̧;���&��[���YN6����i��1�1kޫ�,>��O09��n+�W�F����9�1�֯?e�#3��_ch����V�2��w����~����K0�VDN��8j0�$�\~ �E�f�'
�wn�qDȧ��t����(�/^6�mG�I�RMw%�/X�g��@]=��$��[z�4��C�A��VB��S���t�j�
�� �ѱö��3��)�!t,~ܜH�?���J�J>������f3�4�u�5�߻�M�Z����Ö�Ba��m1���(I'{)�?��GD�/8;C-�Ǆ�]�2߀Ό:5�#^��s3Q\1�!ˁ�m8�P������{�	뼭��Nձ0�'���5}� ;jY��}�D-n��,��9w�IxĎ�;S���h1�ڍ��R�2��'CH?��@��/gﯨ�z����p�j��Sq[Y�pFVԔ�x��n��e����أa؂�IUd.Zl�_����}F�k�� �޹UhH��A��<Ux��_�a�*�΃V}�o���ϝ���r�Ucc�}l�\�z2��A._�������{ߎs�t�ĩS.�*a����1��G��W�%�A*T�=p�1:\���f�����:ީ��½��9�@����c�+���Ü��L��:&TUiX�E�˄9ܱ� ��o;�$��l�Fwvi�h����l���	F14剖�Vb=�5��q��H��ҝ=씩	f��)" �d=Ӂ�?�l((D->qb2��h�]�?�%�B=�cg�!����_���"��Kn8��~��Ci��N���n* ��L����Q��[�!o�{�0�d�f4�)��oYW�5z�!�4�����\?=�~zŪ[����0aKC҈}sTtBG
�؃
��u?a`�	E��6�X��<<O:�X[H�7��W�{�ԕ@�����ߛ|�2�K�P	0Lh��-���uC�t	dC�MO骻����ߌbV���El�v��6�S��E�>�E�u���@=�J��ݨ@C�+��g��TφQ���@=.�D�ۻZ�#!z�VLNڷ	��^���=�s3� ��惬�BrCj��U�0���D�o�����7��Kso�
�f�NH��ߛ�Q�jY� ��ZI���A���\?�����OVS� ���w�6�j<��U=bv4���ܰJ1��/ʁwR���	Ym��kk-�6A����!�><�A�8���v�(�I��vyk"H���,lg�8�P�)�c=:�H��:�� �ĭ�/	�g';�.��d:6xs���>n�Q����ڭ����Ѷ���|�-/	�*��rfL���+�0�� Qb�n��boa��,��'n�
�DJ�r%��i�LKct��?�ܭ9`�2ڜ��2�_=ڨN���}�Ʊd������a^����C�^M���6��zu��I#q
�J'���Kn|�Ȟ������Z���Enˎ) ٪M�4����g�H�� ��bdM�NW�(�8�}1$ɘ%�/#Կc��?+��QFюHk��b��	��Md�@�,�V����ڎ��2�e:���4��<�zTM"�z��#���gKb_ʿV���]P��!��$k$��XJk���߈5W���%V8��4��A�m��X�;�D]#K-��Qa	>����~��J�o☂��L'�	Q�*�0
B��n#��<ʗ\�F"�@
oR�㼯����BJ0?�$�wZ<S+�@HfȊ`T媴���k3B�I�n1B��$�Ě�Ơ�������.�{�����g�����f�m�7�3e��8;���}4V푯/��I_7Kt�	�A���ʼ H���� �!`��#���̍Wh�H<�@"^iiai�?Ț����B� ��O-S��?^.F�"��k�H�S��R�00�;Mo�/v��%m����zﶿH;Jd-��a��j��$[�a�����^�}�0Q�M�Y`�C�Vkfx<��x�%49���b��9��O�V�!�k�\����L?R��B&�	�}�D���>X
��l;�Vd��V��an�yP����v��T��t�0C�Ge� YʋN�Cx5W�p�/�E�&U�dCS��\)>�xw={�W:H
�Qmba�j� ����ٓ��^?
J�6dɀ�x�s��T-v���,-P�{͛����K�f�����4&+�At"6����BaW�f���7��	P6�)��'�\� �/XW���6�����{�6���d�\�pc���@Q�E��Id+����[ �SoΟ�HF�j��uK�]+<�nWs��IߊRMn<ơD�n5�E�o��b!�5��e�_���
d�)dV-}oc��������~��sWyZ�����G��t���ǚ~����}�*���d�"3b���bl����'`�r%�á�3���@~�ɴ�+�^�i�I!e'27U%�e���ln�zr�K�> �^��"��}����B�����1N62�	�A����r��8}���W%	e�
���(u=g���ܟ�tλ��7?����3��4��'3��5\�`�l�!�l/\Ls�m������o3B�K.���f���r�)؜gY�K�:�e`jM'�6�oMz�mf�������2N�f@]}��{�j��H�XNAO&{�X��np�d�L�7	�ý�K�<��zM�Հ[濶.��ά���A8�_y@U`Է�Kd��޴r��H��.� �`�N����<�,��kWN��8 ���b&6�[�z���"npa�)����r�J�B�f�ɶt��������$�.a���߂�����Յ�@�G���.1��n��>nd���h�9ъ�0�I�W�kʹ�7_�<r
�-�L�ַw������O�㵨�<��_���w7"��elj�_�[�T?� I�	�m_�͸b��%����kO(�ضZ*%j2�����hUY��et�x�ǧ\��/������gb�2t�<��;��'���Jb��� �o>f�����7)fwc-yOT0%1O��|M1��XTu�2S,��c�@wK�3v�����C^�Y�A	8c|�����n�B��1�D�5_�IG4��4���C�֩ĨS7iU�f�.�w�����\�s:p0˼s�m?o��B�èԃ�ҟ޻�����(�[��u�X�g���NoiX���9�Q& `D���~Y1�x@��,a�������=;Zt���+;ÇU���I�]҂�P�^NZ�!"�Y���}6�K�?�饄��Q�p���Ⱦ�u��g�՟�^Z����FϽ4�?=�^0;J���%gN�>o�l��y�8j/L��$§�owǔ��c?��8 ��%L<�,�2���^(���랗�i8 �D����i��a�h��*h:=����rHЉz}c��*D�~g`vF-t��h:�!T�+�l��Hzr$�>�hh%Ď_%��YN���{x�CU�NO(.��ɽ��oŕ5�B��b�*��&�C���#3��R[��&�㦗�^��>�[���*AW����Ebn.��	'���vY�!�n�]�t�v���a�~��ʠ��������p,4jѹ�z������͟��ܪ�������g�oE6R3o�A�@���SY����($�m�Ojc�r���9;5�s�ͣu��U���k�x�I��}H��yi�kɝ�$�D�;',� VK��:�*)W��k��1^!u��. �^�<�	��ٶ���.<��DXYk���+�3u�"Z'�}a�3E?'���c-��� J����bz�䤮�����éE\���3&��N�0��&�6���N@�Ie6%_4�0��D{�k?�����\d#�d�zX�K~�e��x�3W��]���ř,\Z�42[�1����9�A<���<������G�%^W�N>H�gtR�~u�K����Z��
�:Nh��k� ��T�*�c������D����`cǏ�3�����XQ�9�l9��>$4	&.p,�eё�%��"�j��<�w��E�S$+8�{)鲠
��]�f&�O��-�l5^��&y�I��6�hi��Ҕ��ͅ�XGڀ@&�6W�߃&�˕2psA�9��Yp�eC��\���>y�WCiz/��d�-��ћ��1�ښ[�+����c�x`+Sr�FDh%d�;=���T�/F:e�gO�B�ρ�7p���ٴ54�-52��Y6�\�K
1M<���}M��e)l���&�o��K�B�RIgZ�������h�-h\5�ܓ���lh6v{�Mk���X0:Jü(�Hg i�_�̝Y;IC?!��}�T5N��Q{��<�>�� ��@����d O�a����#����AV��5�6�}��>��E�-���7�&��8\Os�E:��S��9�*Ad,�X�LO���x�����|�i����q;5�l�&L{�d8�����^�mC]���5D�:���������#<��"�C��2g{gkk��cp2�`�vAvf��uY��%Q ��1�U~)��:6��G��:�I`4 L��9��U�ClK�<l+�V܊u*/J���li���߀�{y�n1O�4 ��t�Qv�(2�_�j�n�.�L~�r��'������A�
��o�W�_=t�Wx���_��P�Ɂ��e�b�>����"��;x�&��>�ȼz��;ce.���5�es�0�❢��4qI���-Z��W�F<���}�A*���=�M.XBز,U&l�]C,]x��$U�{�"VBd�=.���#�wEW&��%<2!��K�3�߱��}ħ��������;�dj���f#S#�^�Q22�ZC������\]�0f��4c�OMMV�b���2dXlxVHYEB    fa00     cf0!8F�����u���SH+���Xox���7�q]�uq�p��mT��d�_�U����ݱ�����x{�Jq�2G����	�-p�
�j7aLX$<�u7xW3[]�w��Qj�?]aI�\��s*�8���I��X����C���t���|՝<E��Q0:���
��᲻W�U$��Vb2p����%G�j,����
����t�ͼ`˄w��.�r��u��ch�%xE�Ѱ���ؽnj|䙋�ï��������ס�R��g�����T;�&=EFy�*/-=h� 7b���Ri(f��
_��$�>��%�
s{z��TW�7�[��	�A�zƈ~��w�+����Ae����<$���qX��b�l�\��Ore@�(�͕�4����)��kx�g����nZ�4�V� �B�f�\�,���(�YG�mE��t���s�@���-����<K=F�CjY�.#	��&�b�g�M!�#�HMR�5%��������ƪ��֣MK�p}�x���^�F����ۧ/Ƴ�l�>n�k��h��t�'XQ���T"O#s�����Pz��Qk
��_Y0�xw?�Fag95�E��y��x&��jf`��S�e��E,���J������-�<5�u�����cnoh����vʹsQ�;�*Ϲ�~�O�wu`a��t��PhD���uz,M�Q���7�*,�)�u��I�f�DP��o�/
o�[�?�Zӌ�מ�?��F�2f� �� �[��篁Y��ڬ��(A�'`Ef���Q�K	@9��z t�t��<e��2�c�>�?x�t�B���܅@ԯ�����@��D�F���.��:���y�Q�x?�rWpmY���ޞQp�g8b3����B���sQ}q��SH�$y����%��C�'���1�.S{�����Y�����~�PYR31{K�ъ`·���M���w��<��\��lȶ~�}'M:|b�;���B��t���f��5�	��)���D�0�����O<���>n%�t"���]��[!���n��Y���4z�>��,��y�����d��ލ�U��}i�ڭ0����
���a��%E&>���3�u/����w6�j �\C��K��;�y@���c����@����Q,�/��z�(5�n���j��X a�M�eȌsGG�`S(�<��
��V����Tc��]�	�=��x�^b��C��<N`E���_~؛�#ϝ��I�'��n���L�k�pXm�T���%���2�VN�iq^���IB��Q��׈Ԕ{�?4����F�s�8>U���n�k��9�1/LO8���0`w�O�PjiТ�X(�
�@�߷�}�J��;��X����wt�;��%��zc��jسz腆BG0��. �M��;��x@@�4��2�Ty��끄���/ *r��O��`��/7�PO�n��T�7YP�/�k)�3�}�~�c
�WL�Gy�%2`^�Y�����Kg�!ǳ��s����'�� 8C�cM`6�JQ�}�1�1ˑ,A�g6�[�p��qYk�޸�J؟LyO���α��6�-fivr���6{Ҟzà^p�Kj�A%�����bv"��d���f����Dd{¥k��>�4� ��i}�g�}����=t�;�1�ھ֦õE@��S����`�~�aP2��0-���,�5x�D�?ٱ#�[F��9���s��c7��g8D@l�G�?�E��t^��[.�����̌�L� ����Q�������8s��}u�\�;��/�	| gf�����JeZ:�2�%l�����گ���}-t�����@�!J�x�%UF����zm_AX4[V��)ȽTT�Y�:5q�d�f�B-2h�5l&��>N���!y�wN��I�*c�'�?<�z+��(0��+a	�����s�#�]G��و7��Wg $̖}Ӟ�l�u�<�����z{����D"tY�r^�A ��ul#�{��~��3��?���<�B���!���M���
{(�Y�B�OJ]2M������B��C�yh��+���(&t)���-J�*FW�=~����Ĵc-�m�qD%�jM�d�g�>���?�I�RYp�>�-�k�(E�7�9��č��]��)��rWk�OaV��{. $[�aq�At��"UPA����꟧%�֧�1L3��Ov@��������E�Xd�_��Z�-F6c�(ԋ��e�jbv��s s���մ��bP�?�n7y��WDK�8cr�W'|�?�W��!��0���V)KgV��&��"6�;?N?5tW�	�S�z��5��
M�{b��+*ѹcO�ͳ�N]n��;h�f�6U�~���Fx���ŷ��������c'��S��E��4N�B���x��m�mB��K��ʆ�G�d���jV-s���J�N�z�
�yd����T"SI�hu;J/_�<zgZ$��g�@zóQXu�K�lh��=|6/��{u��YhA��s�wm��=P���{�<��u&ѧl�e�`��P��a��������oRK\���)�C23GN�}b���iZC4�QP�؉�ۖR��+���L?g5P#1ߒz3E���6���ԗ�ShT2�*t��⼣d�gP��r?�!��v"�0��U(�0�׼V���AE���g�K�j�$��1�e��~��G9<�c���l�����Ǘ7��F\#�ӝ:���_D}�5d\�+_�kA��?�E
Y�$7e����y�n�h���J1��82�(1��Ѵ������b���q�߳�m��Y��Y��fK�iAF�㶍��JFF5�W���x#�$9FD��@���K��jeT��
�����-�2�����!S�'��7K4��#��j���sy(5�*o&B����Si7��'�Hi�TBJ���W�M�&���Tp��uv'yj�h�GNgű�|��DG�+�$�ж0ѕ�:��ʪǤO��Vk�h(V���t���Ck�l4�҇�ਖ਼ 5D������?�^P%�
�޼J��N 3K�A�AcT��V�����Y��pc�gK����hP��
��q3Jp��|���)x�s��O�7&��-�r/��[6�:Ng�8T��\�Ew}��K'��ӉN�8���r���

E�Y�)��!�ۛcr��I�!=A�)T´�˚ڤ��Q@�_{"2��AR_��J�F^ǩИf聤p������.m]:���,Oʲg��􀯄���R1s�COF]���p
Ucm3 h��Z����n�\�)�*n*XlxVHYEB    3981     4d0Q�曛����3�J���}��I��緙� E>��8�6�v��Z��mJ�W�){���z}��'��D{�������EgAG�^��(�����e�5z�a����2��}�u��Ү�Y,h5GQ3�����2��.� ������y�2V4x���W�/ǋ�m�a�d���9Q���|v߸�9ξrK6�(�:۶&:b��cBq�m�-Fjb	���T�I�#10M����JKU�,�-V���CL�t�>��I&��R~�4�W(�r	�-m�e2�8�_�����+�D�.4�J�Q�V�s5}L�@qy}ze,���M������|�h� �o�#A��~����`�9��~{����n��]���i�<��:�{EH�(af�?��\T����������si�ϓ�K*BCWwH�\�L!h��%5 ��
�F ���Z�%Y���+�#�0l�E&IU�ۮ
�z��Jd�,��1�>��bf�LW/��TZ`�p�����(�t����Z�� ���z|�`߽d�:� �68��)�!�P̀�-��{G/]�4trezw���S�^o����ﮜ?�L��E�`FQ�÷9zm�������5b�l����$C߯�a�x!s���*މ���Y������0P�J������d��'Jd��=aDƊ�w��o�*
��^�2dD�mwJE
{�x'�$-�5��P��	|��v+b��x�ӧ�Zz�ۮ���E-ʜ26� 0X���9�شe�P�m�5E��F<c���g<⟊8�a;��$S�?>�#"�%���W��,���vd���������'-[^d���Ak���<��y7���I�������VM���1X�,��DuYe?G1 ��tOES�Cl~��l>�;�.��v�F#H��6B���<�\��tY��<����RM04��>ol���H�~zf#� �d����Q�'x+�-�А�f�D��K�^�_�ݏ *��^\����-g��yUtYx1�O�����v^�7,H�Ds<��+��	
K\g�L�O�y��MF�A��[�h�ˍ�ߠ�!�R0 yX��Mm��#
e����n,!����ο-���;���0�C��6��r }��C5]ּ�|D�X~�>6B���~lԘ�gm�⎹�6�����1q	+7��M	;��<Q?�G|��C� �.\�I��0�����l�4�����lfk��
%ޗq: