XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���ߟ�
+u��+Dwӭ���H_p�wGǔ��I�b���5t���餮Z�C�U�&'�b��REh��{�"c.�� ;���ئ�lA�C� �B�8�f��E�Lp�����.�ԲN-ނN^���(λ/vv3Ɵ�����bS���d�@��V��+��y�qOf-ю�ߧ6��Vy/�qR�4!|���iL�'��3){AR,j�z.�^TX��)ܓ��[Ǩ�����igs.tK�k���w���!O~�o惚j~T8� >������-���z�}�8���E��;�,� �f�ґ�Ogv:�+��_���OR#-x�.}U��l����]S��q���-�M��<O��%3���Ąl�Vt���� e��	|�_<�{dڱ��³x�Դ�%��	źUe�3�~qe��9�iq��=����I�GS��T&���ā1�(30�mum,I�/կp��;��9�o��8^�!�l*���a��))5I�$�
�´������jxe�� �C �B�>�f����r,s�������^'��j��ӂޒ���i��r��y��87n�}i6a�(�6XŒ��~�Nָ�O! �#�`:�R%�=�@>v�ttg��/o������5/ZW<b��)a�:MO��~t����`�39-��F�cmK-/�0��0(�y<r��9oʘt3!��vo�ƨi����qC1Q��9����ˊ֨G�LO��ł��|mL�ă�̕�K�pp��1�ӳ���1�W0�(C���#W�\�[2XlxVHYEB    5b76    12f0�&���jA�<�uMO�ﴕ���+�xR�.�u�~����cF{���w����6Wߨ%�M�k�Ъ�n<�{˕��+����#��0�e�����N<���<�E���8���Ӂ'����ȡ#[T�D��������G��MŴȮK��5�ޜw��cHx�O`�;J�(��R�T�"ID�g��a�p8o�˗.�h��,W�m�vw�6b�l)w�do���?��o��UqG�>�sgw�)�7?��vIH�8HU6V��*X*���j<\�}I��OI��j*P����i^L�6�,�n`�W<�u]�M�g��E1j6fbE�)I�o��<��u��-�K'�r���QG�6&�jg��$6���ex3�}5z:���T�D�]!B.X~�&̒"�9~ܬqcRļ�(�(���4�Q�8�o�%c �[��×sa�o)T���4���$�\�?��$"��9��a��W�� ��6�g� �ʓ��F8Y2<��<�'Gx��//��:&��+�J�D���#v��2�����x����������ĐI[�T:<p�=q���ڵ�-00K��{�4�z�����h~)Ds��S4�Т�������l�;{���W�yhb�b���fD���h�x3�@3���`�'c2����f�r�s޼��#�r��+s��0sb�:���=&W��E��|>OE��a�����b��R��{m��r�0��ge+��)� �]�Qf���~k:q��R~J�}%ne蚖]. ��K�G�YaƟH=���э����ь���%RSkvk�6�;iS����'�w���?qm��5�[_��2C���갰��oW-��_Ҝ�K�	����o9Љba���n�&�k�6h+C�W4
�l<HW{��/�����R��^���Q���b?��|��q	@K�n�&���b2�UQ����6/1��I��AN�1E��nL��c,��N���Jw�a��S�,�rr����z@E��5��y�5RM?���~��j�d��j��T��u�r��k�ڢ�g[����F��%N-�����b�W]g��?8;��Zv��ǅ'4c��y]��XG@��=�g���s���=�W�N|"�b���& ����#�A���~: ��w�|��:1����4�����[��E=������Cw�𧎵8I���7zצ�x�g��  ��̝��H������Y�!�\������ɠ�-�Z�����K$��N*�C���4�B�&�ʛQ�D�) .�f�������ь�S��U���D����C��M��Ƨf����vN�Y�%M������X�J5Ѯ<�k�Ao��2��[�l>і���+JSZ��Z7�H��+�>Q1`��)�<R=��.Uf���JvQD������b's�GX��Zw�SaF�&6��bD3[��To2�A)���;��P��E5u֑��{* �����Z����SST~)��'Tԗ�*t��9�i|"�\��Fj����m��ܹ��P�X�w��#�%����F��U w�r�'��[Nk���
vƁ���73�s��5N2��G��hѶ���y��K%������$=�kЊ�m�J=�
��q��Y��� ~�	6��?��Q�[��q������^O���8�r�H0Ȣ���<.n��;�V��+v��":�����C
�6���ZX�˙�Ug���`��e(�E�+vzX���K��z�l�@��-R-���3/�@�_������>+��f��X�֏o
��D�vr�]>f��&�1�p"8v��u.�lP�����>�u�j�y�w���?�fb=�����<�P��L�9�U�?���)�I�r��=������S�<OP�,��%��7�5���� ��'��*�|�]yGgz���h�w7j�"�-N��sD˪��Yfrg9�-\��V���|�PǾ�pc���\����~��b�4�_�`�/�k"Z�N&=����+~��L˲������O��_�8�T̒����OF)79�_tߋ���^�c��5�@馰а����S'�z�^��EF\A5��'ʡ��3P1Cw�.������</�xU0�L���a��&�+��08��t��qJ=ݗ�ږݶ��<��*eŕ�����͓�۱�u��o�ɿ��:J04��R:o��x�i���&(*g	
����9h	��+ލ�6k�ۡ��H�}Z$�XI���� ?2	�X~�?�*�ʷ���>�O�����H�4s�y@��2���vu�9Cn���?�]")�Hy�;q� ��ut�W��U��My�9bG��>Թ<��`���H/a��7fNL��iUX��yG-���� ��a��k�e�&���@�(h��
'�$�P7���'�>)��a4�^�e2y�L⺓�v-X�u���G��
|zR��Z�ٴ��'�MN?�443�t���6��HQ�݄�jqu�K�<�e�Z'ˢO%�=bn��}u�c��&O[�&�4��r}l�ە `�E�p� �5�\��2o
���뱆�~̐�5k��I5����=1N��/Y���#y�M۩Q��[�6Hx8 �*�v����k�u��hf+�L�+-U���[�R��R|�H̟��o��y���ɡ|Ql�zh��a��~�y�)�ҭr��M���@�q�I�/:]�#��|A��N���X�!��jr3��探�WAR��.�
��FpGaG��,�@���RbI�o���Fǔ����<�9�G7[lU���L�c�8M3�z��[�[:i�PwTd�ڵ��²�
-������m1��������Uj2	T>HҴcM��a���I���O
�C���O¤��d��VZ�}��i�x�.���<2�T�;��AA�F���^�	���led��n�ό�� {��1�G]����1�֛*Ko@�I\T;��'�������LZN-)�Q�P��pqr��
�?�WtS-8�_o"cu�՘	�Vp[*Z�Y�ic�����C�3���g�˱�R���Ϥ�Z��Y���w��P����m#��?��mbƜ$����e�i8>���o9ގ�PQk���;':��Dc��wf}z��(@v�i��G�c���9X�u�Lsu�
��O/F�ΩQCC�H�p�g��Ջ�P��gP�=QW���k��x�XitR���ثM��=���(R��j�(�g$�3�k���m�%�Q��7a60��E�Y���R4ߚs���y_q��N�s���r��i��Qܸˀs�	�4�P,���H�8���!6��:_�Oc�NX���=��$�!�ZE��0|oT����-��ՔX;�Uh�0��P�T>온�0�]rN&��B�q��S���+��_�EA��*��a�GtN��L���� _�
a�}@��p�W�:a�yPu�����KOՔ�Ro�b������"@*������<�z�%3޳_Ď�6X��޹�oF>�G��8��6�<��pd��������9����T'1{��D��B�F�f�r���Iժ@�[��Ls��l�8&� �3��3�P��N_�5|��Ӈb��e�����n�Yvm@��>X%�� ĦJoa܋��j8���]m)N�=k.9��r��J�� =zo_$k���
FEB&��O��Yey��JW3-*���Eԟf�[rY����.���$t'�LřW17#�p|!�)�F��n��j6i9����A��+�p$���B<�l�c�Җ���� ���O�\PGK�(��/[��eT��2�6`ewq]�94��w�4�����a�a^�8z�
��aDxj��ŏG�S��3ÿ;�F��)�]��qt<����}��?L��f�^�R�v"H�4t��H���1��՚2Z��^R�me�R݅6�]��Y<�U�D>��ś�3ޚ�q�1�D0�r�*��-XNP���T�����Dk�\o�p��K���?�V�`�L�yy\���5;H�-4�7�8m$y����~#'$5���p/�?qP ��J�,��O6YD�`��E�w:�Kz�|�)������0�yJNؗo=���V������O/��?=����.�zk2���bCv2J�]<��]$�q��t�'��A�x��C�2��j��(q�K.Z{!�!�ט)��6(�cD�o�l�ò�U�:{�]���z�-��)Ě�tʛ�����
�P_!c} �����-�`9��L��%�"��WOL��Xy�]#mk���Ԩ;Qfa�� ���ÉmC�O)��}�� z����3�@����4����.���JIv��d���(�wc�3z���#C�|'�{�f���f���eW%7��)�t�ƿLC�5c�;g��ֲ� ��p�#ݗ��+\/��̊@%<�T�j��� &%;}2w�LFB�U������fc���rN���*˺��ӷ �xX����M8F�1f�'T�%��qۤN'L
��ծ��S1�;����U�?���P7�V�rH��8.[)�'n����(���4��e�����N�h�����-���ʸ�@�&�����1�h�8����U�eD�V�.�����w�Wb�T�p}>R,�::wl��7��b8�3����{�R��Vd=(e�ݙ�[J�N)���!�{���$�F��H<T���tf�V���i���@�\7K��2+��`f�s�@/ c��xJaFfCo�.�c��Hi�7S�}zi)�]�-C0���Eh���6��:Q#;kEd!��r�Ғ@�:SB:�����L9�,J6gO�w�M��